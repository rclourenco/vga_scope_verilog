module WaveRomTwo(
	input wire [9:0] address,
	output reg [8:0] data
	);

always @(address)
begin
    case (address)
        0: data = 9'h0FF;
        1: data = 9'h116;
        2: data = 9'h12D;
        3: data = 9'h144;
        4: data = 9'h15A;
        5: data = 9'h16F;
        6: data = 9'h183;
        7: data = 9'h195;
        8: data = 9'h1A6;
        9: data = 9'h1B5;
       10: data = 9'h1C3;
       11: data = 9'h1CF;
       12: data = 9'h1D8;
       13: data = 9'h1E0;
       14: data = 9'h1E7;
       15: data = 9'h1EB;
       16: data = 9'h1ED;
       17: data = 9'h1EE;
       18: data = 9'h1EE;
       19: data = 9'h1EC;
       20: data = 9'h1E8;
       21: data = 9'h1E4;
       22: data = 9'h1DF;
       23: data = 9'h1D9;
       24: data = 9'h1D3;
       25: data = 9'h1CC;
       26: data = 9'h1C5;
       27: data = 9'h1BF;
       28: data = 9'h1B8;
       29: data = 9'h1B2;
       30: data = 9'h1AC;
       31: data = 9'h1A7;
       32: data = 9'h1A3;
       33: data = 9'h19F;
       34: data = 9'h19C;
       35: data = 9'h19A;
       36: data = 9'h198;
       37: data = 9'h197;
       38: data = 9'h197;
       39: data = 9'h197;
       40: data = 9'h198;
       41: data = 9'h199;
       42: data = 9'h19B;
       43: data = 9'h19D;
       44: data = 9'h19F;
       45: data = 9'h1A1;
       46: data = 9'h1A2;
       47: data = 9'h1A4;
       48: data = 9'h1A6;
       49: data = 9'h1A7;
       50: data = 9'h1A8;
       51: data = 9'h1A8;
       52: data = 9'h1A8;
       53: data = 9'h1A7;
       54: data = 9'h1A6;
       55: data = 9'h1A4;
       56: data = 9'h1A2;
       57: data = 9'h1A0;
       58: data = 9'h19D;
       59: data = 9'h19A;
       60: data = 9'h197;
       61: data = 9'h193;
       62: data = 9'h18F;
       63: data = 9'h18C;
       64: data = 9'h188;
       65: data = 9'h184;
       66: data = 9'h181;
       67: data = 9'h17E;
       68: data = 9'h17B;
       69: data = 9'h179;
       70: data = 9'h176;
       71: data = 9'h175;
       72: data = 9'h173;
       73: data = 9'h172;
       74: data = 9'h171;
       75: data = 9'h171;
       76: data = 9'h171;
       77: data = 9'h171;
       78: data = 9'h171;
       79: data = 9'h172;
       80: data = 9'h172;
       81: data = 9'h173;
       82: data = 9'h174;
       83: data = 9'h174;
       84: data = 9'h175;
       85: data = 9'h175;
       86: data = 9'h175;
       87: data = 9'h174;
       88: data = 9'h174;
       89: data = 9'h173;
       90: data = 9'h172;
       91: data = 9'h170;
       92: data = 9'h16E;
       93: data = 9'h16C;
       94: data = 9'h16A;
       95: data = 9'h167;
       96: data = 9'h165;
       97: data = 9'h162;
       98: data = 9'h15F;
       99: data = 9'h15C;
      100: data = 9'h159;
      101: data = 9'h156;
      102: data = 9'h153;
      103: data = 9'h151;
      104: data = 9'h14E;
      105: data = 9'h14C;
      106: data = 9'h14A;
      107: data = 9'h149;
      108: data = 9'h147;
      109: data = 9'h146;
      110: data = 9'h145;
      111: data = 9'h145;
      112: data = 9'h144;
      113: data = 9'h144;
      114: data = 9'h144;
      115: data = 9'h144;
      116: data = 9'h144;
      117: data = 9'h145;
      118: data = 9'h145;
      119: data = 9'h145;
      120: data = 9'h145;
      121: data = 9'h145;
      122: data = 9'h144;
      123: data = 9'h144;
      124: data = 9'h143;
      125: data = 9'h142;
      126: data = 9'h141;
      127: data = 9'h13F;
      128: data = 9'h13E;
      129: data = 9'h13C;
      130: data = 9'h13A;
      131: data = 9'h137;
      132: data = 9'h135;
      133: data = 9'h132;
      134: data = 9'h12F;
      135: data = 9'h12D;
      136: data = 9'h12A;
      137: data = 9'h128;
      138: data = 9'h125;
      139: data = 9'h123;
      140: data = 9'h120;
      141: data = 9'h11E;
      142: data = 9'h11D;
      143: data = 9'h11B;
      144: data = 9'h11A;
      145: data = 9'h118;
      146: data = 9'h118;
      147: data = 9'h117;
      148: data = 9'h116;
      149: data = 9'h116;
      150: data = 9'h116;
      151: data = 9'h116;
      152: data = 9'h116;
      153: data = 9'h116;
      154: data = 9'h116;
      155: data = 9'h116;
      156: data = 9'h116;
      157: data = 9'h115;
      158: data = 9'h115;
      159: data = 9'h114;
      160: data = 9'h114;
      161: data = 9'h113;
      162: data = 9'h111;
      163: data = 9'h110;
      164: data = 9'h10E;
      165: data = 9'h10C;
      166: data = 9'h10A;
      167: data = 9'h108;
      168: data = 9'h105;
      169: data = 9'h103;
      170: data = 9'h100;
      171: data = 9'h0FE;
      172: data = 9'h0FB;
      173: data = 9'h0F8;
      174: data = 9'h0F6;
      175: data = 9'h0F4;
      176: data = 9'h0F2;
      177: data = 9'h0F0;
      178: data = 9'h0EE;
      179: data = 9'h0EC;
      180: data = 9'h0EB;
      181: data = 9'h0EA;
      182: data = 9'h0E9;
      183: data = 9'h0E8;
      184: data = 9'h0E8;
      185: data = 9'h0E7;
      186: data = 9'h0E7;
      187: data = 9'h0E7;
      188: data = 9'h0E7;
      189: data = 9'h0E7;
      190: data = 9'h0E7;
      191: data = 9'h0E7;
      192: data = 9'h0E7;
      193: data = 9'h0E7;
      194: data = 9'h0E6;
      195: data = 9'h0E6;
      196: data = 9'h0E5;
      197: data = 9'h0E4;
      198: data = 9'h0E3;
      199: data = 9'h0E1;
      200: data = 9'h0DF;
      201: data = 9'h0DD;
      202: data = 9'h0DB;
      203: data = 9'h0D9;
      204: data = 9'h0D6;
      205: data = 9'h0D4;
      206: data = 9'h0D1;
      207: data = 9'h0CE;
      208: data = 9'h0CC;
      209: data = 9'h0C9;
      210: data = 9'h0C7;
      211: data = 9'h0C4;
      212: data = 9'h0C2;
      213: data = 9'h0C0;
      214: data = 9'h0BE;
      215: data = 9'h0BD;
      216: data = 9'h0BB;
      217: data = 9'h0BA;
      218: data = 9'h0B9;
      219: data = 9'h0B9;
      220: data = 9'h0B8;
      221: data = 9'h0B8;
      222: data = 9'h0B8;
      223: data = 9'h0B8;
      224: data = 9'h0B8;
      225: data = 9'h0B9;
      226: data = 9'h0B9;
      227: data = 9'h0B9;
      228: data = 9'h0B9;
      229: data = 9'h0B9;
      230: data = 9'h0B8;
      231: data = 9'h0B8;
      232: data = 9'h0B7;
      233: data = 9'h0B6;
      234: data = 9'h0B5;
      235: data = 9'h0B3;
      236: data = 9'h0B1;
      237: data = 9'h0AF;
      238: data = 9'h0AD;
      239: data = 9'h0AA;
      240: data = 9'h0A8;
      241: data = 9'h0A5;
      242: data = 9'h0A2;
      243: data = 9'h09F;
      244: data = 9'h09C;
      245: data = 9'h099;
      246: data = 9'h096;
      247: data = 9'h094;
      248: data = 9'h091;
      249: data = 9'h08F;
      250: data = 9'h08D;
      251: data = 9'h08C;
      252: data = 9'h08A;
      253: data = 9'h089;
      254: data = 9'h089;
      255: data = 9'h088;
      256: data = 9'h088;
      257: data = 9'h088;
      258: data = 9'h089;
      259: data = 9'h089;
      260: data = 9'h08A;
      261: data = 9'h08A;
      262: data = 9'h08B;
      263: data = 9'h08B;
      264: data = 9'h08C;
      265: data = 9'h08C;
      266: data = 9'h08C;
      267: data = 9'h08C;
      268: data = 9'h08B;
      269: data = 9'h08A;
      270: data = 9'h089;
      271: data = 9'h087;
      272: data = 9'h085;
      273: data = 9'h083;
      274: data = 9'h080;
      275: data = 9'h07D;
      276: data = 9'h07A;
      277: data = 9'h076;
      278: data = 9'h073;
      279: data = 9'h06F;
      280: data = 9'h06B;
      281: data = 9'h068;
      282: data = 9'h064;
      283: data = 9'h061;
      284: data = 9'h05E;
      285: data = 9'h05B;
      286: data = 9'h059;
      287: data = 9'h057;
      288: data = 9'h056;
      289: data = 9'h055;
      290: data = 9'h055;
      291: data = 9'h055;
      292: data = 9'h056;
      293: data = 9'h057;
      294: data = 9'h058;
      295: data = 9'h05A;
      296: data = 9'h05C;
      297: data = 9'h05E;
      298: data = 9'h060;
      299: data = 9'h062;
      300: data = 9'h063;
      301: data = 9'h065;
      302: data = 9'h066;
      303: data = 9'h066;
      304: data = 9'h066;
      305: data = 9'h065;
      306: data = 9'h064;
      307: data = 9'h062;
      308: data = 9'h05F;
      309: data = 9'h05B;
      310: data = 9'h057;
      311: data = 9'h052;
      312: data = 9'h04D;
      313: data = 9'h047;
      314: data = 9'h040;
      315: data = 9'h03A;
      316: data = 9'h033;
      317: data = 9'h02C;
      318: data = 9'h026;
      319: data = 9'h020;
      320: data = 9'h01B;
      321: data = 9'h016;
      322: data = 9'h012;
      323: data = 9'h010;
      324: data = 9'h00F;
      325: data = 9'h00F;
      326: data = 9'h011;
      327: data = 9'h015;
      328: data = 9'h01A;
      329: data = 9'h022;
      330: data = 9'h02B;
      331: data = 9'h036;
      332: data = 9'h043;
      333: data = 9'h052;
      334: data = 9'h062;
      335: data = 9'h074;
      336: data = 9'h088;
      337: data = 9'h09C;
      338: data = 9'h0B2;
      339: data = 9'h0C8;
      340: data = 9'h0DF;
      341: data = 9'h0F7;
      342: data = 9'h10E;
      343: data = 9'h125;
      344: data = 9'h13C;
      345: data = 9'h153;
      346: data = 9'h168;
      347: data = 9'h17C;
      348: data = 9'h18F;
      349: data = 9'h1A1;
      350: data = 9'h1B0;
      351: data = 9'h1BF;
      352: data = 9'h1CB;
      353: data = 9'h1D5;
      354: data = 9'h1DE;
      355: data = 9'h1E5;
      356: data = 9'h1EA;
      357: data = 9'h1ED;
      358: data = 9'h1EE;
      359: data = 9'h1EE;
      360: data = 9'h1EC;
      361: data = 9'h1EA;
      362: data = 9'h1E6;
      363: data = 9'h1E1;
      364: data = 9'h1DB;
      365: data = 9'h1D5;
      366: data = 9'h1CE;
      367: data = 9'h1C8;
      368: data = 9'h1C1;
      369: data = 9'h1BA;
      370: data = 9'h1B4;
      371: data = 9'h1AE;
      372: data = 9'h1A9;
      373: data = 9'h1A4;
      374: data = 9'h1A0;
      375: data = 9'h19D;
      376: data = 9'h19A;
      377: data = 9'h199;
      378: data = 9'h197;
      379: data = 9'h197;
      380: data = 9'h197;
      381: data = 9'h198;
      382: data = 9'h199;
      383: data = 9'h19A;
      384: data = 9'h19C;
      385: data = 9'h19E;
      386: data = 9'h1A0;
      387: data = 9'h1A2;
      388: data = 9'h1A4;
      389: data = 9'h1A5;
      390: data = 9'h1A6;
      391: data = 9'h1A7;
      392: data = 9'h1A8;
      393: data = 9'h1A8;
      394: data = 9'h1A7;
      395: data = 9'h1A6;
      396: data = 9'h1A5;
      397: data = 9'h1A3;
      398: data = 9'h1A1;
      399: data = 9'h19E;
      400: data = 9'h19B;
      401: data = 9'h198;
      402: data = 9'h194;
      403: data = 9'h191;
      404: data = 9'h18D;
      405: data = 9'h189;
      406: data = 9'h186;
      407: data = 9'h182;
      408: data = 9'h17F;
      409: data = 9'h17C;
      410: data = 9'h179;
      411: data = 9'h177;
      412: data = 9'h175;
      413: data = 9'h174;
      414: data = 9'h172;
      415: data = 9'h172;
      416: data = 9'h171;
      417: data = 9'h171;
      418: data = 9'h171;
      419: data = 9'h171;
      420: data = 9'h172;
      421: data = 9'h172;
      422: data = 9'h173;
      423: data = 9'h174;
      424: data = 9'h174;
      425: data = 9'h174;
      426: data = 9'h175;
      427: data = 9'h175;
      428: data = 9'h175;
      429: data = 9'h174;
      430: data = 9'h173;
      431: data = 9'h172;
      432: data = 9'h171;
      433: data = 9'h16F;
      434: data = 9'h16D;
      435: data = 9'h16B;
      436: data = 9'h168;
      437: data = 9'h166;
      438: data = 9'h163;
      439: data = 9'h160;
      440: data = 9'h15D;
      441: data = 9'h15A;
      442: data = 9'h157;
      443: data = 9'h154;
      444: data = 9'h152;
      445: data = 9'h14F;
      446: data = 9'h14D;
      447: data = 9'h14B;
      448: data = 9'h149;
      449: data = 9'h148;
      450: data = 9'h147;
      451: data = 9'h146;
      452: data = 9'h145;
      453: data = 9'h145;
      454: data = 9'h144;
      455: data = 9'h144;
      456: data = 9'h144;
      457: data = 9'h144;
      458: data = 9'h145;
      459: data = 9'h145;
      460: data = 9'h145;
      461: data = 9'h145;
      462: data = 9'h145;
      463: data = 9'h144;
      464: data = 9'h144;
      465: data = 9'h143;
      466: data = 9'h142;
      467: data = 9'h141;
      468: data = 9'h140;
      469: data = 9'h13E;
      470: data = 9'h13C;
      471: data = 9'h13A;
      472: data = 9'h138;
      473: data = 9'h136;
      474: data = 9'h133;
      475: data = 9'h130;
      476: data = 9'h12E;
      477: data = 9'h12B;
      478: data = 9'h128;
      479: data = 9'h126;
      480: data = 9'h123;
      481: data = 9'h121;
      482: data = 9'h11F;
      483: data = 9'h11D;
      484: data = 9'h11B;
      485: data = 9'h11A;
      486: data = 9'h119;
      487: data = 9'h118;
      488: data = 9'h117;
      489: data = 9'h117;
      490: data = 9'h116;
      491: data = 9'h116;
      492: data = 9'h116;
      493: data = 9'h116;
      494: data = 9'h116;
      495: data = 9'h116;
      496: data = 9'h116;
      497: data = 9'h116;
      498: data = 9'h116;
      499: data = 9'h115;
      500: data = 9'h115;
      501: data = 9'h114;
      502: data = 9'h113;
      503: data = 9'h112;
      504: data = 9'h110;
      505: data = 9'h10F;
      506: data = 9'h10D;
      507: data = 9'h10B;
      508: data = 9'h109;
      509: data = 9'h106;
      510: data = 9'h104;
      511: data = 9'h101;
      512: data = 9'h0FF;
      513: data = 9'h0FC;
      514: data = 9'h0F9;
      515: data = 9'h0F7;
      516: data = 9'h0F4;
      517: data = 9'h0F2;
      518: data = 9'h0F0;
      519: data = 9'h0EE;
      520: data = 9'h0ED;
      521: data = 9'h0EB;
      522: data = 9'h0EA;
      523: data = 9'h0E9;
      524: data = 9'h0E8;
      525: data = 9'h0E8;
      526: data = 9'h0E7;
      527: data = 9'h0E7;
      528: data = 9'h0E7;
      529: data = 9'h0E7;
      530: data = 9'h0E7;
      531: data = 9'h0E7;
      532: data = 9'h0E7;
      533: data = 9'h0E7;
      534: data = 9'h0E7;
      535: data = 9'h0E6;
      536: data = 9'h0E6;
      537: data = 9'h0E5;
      538: data = 9'h0E4;
      539: data = 9'h0E3;
      540: data = 9'h0E2;
      541: data = 9'h0E0;
      542: data = 9'h0DE;
      543: data = 9'h0DC;
      544: data = 9'h0DA;
      545: data = 9'h0D7;
      546: data = 9'h0D5;
      547: data = 9'h0D2;
      548: data = 9'h0CF;
      549: data = 9'h0CD;
      550: data = 9'h0CA;
      551: data = 9'h0C7;
      552: data = 9'h0C5;
      553: data = 9'h0C3;
      554: data = 9'h0C1;
      555: data = 9'h0BF;
      556: data = 9'h0BD;
      557: data = 9'h0BC;
      558: data = 9'h0BB;
      559: data = 9'h0BA;
      560: data = 9'h0B9;
      561: data = 9'h0B9;
      562: data = 9'h0B8;
      563: data = 9'h0B8;
      564: data = 9'h0B8;
      565: data = 9'h0B8;
      566: data = 9'h0B8;
      567: data = 9'h0B9;
      568: data = 9'h0B9;
      569: data = 9'h0B9;
      570: data = 9'h0B9;
      571: data = 9'h0B8;
      572: data = 9'h0B8;
      573: data = 9'h0B7;
      574: data = 9'h0B6;
      575: data = 9'h0B5;
      576: data = 9'h0B4;
      577: data = 9'h0B2;
      578: data = 9'h0B0;
      579: data = 9'h0AE;
      580: data = 9'h0AB;
      581: data = 9'h0A9;
      582: data = 9'h0A6;
      583: data = 9'h0A3;
      584: data = 9'h0A0;
      585: data = 9'h09D;
      586: data = 9'h09A;
      587: data = 9'h097;
      588: data = 9'h095;
      589: data = 9'h092;
      590: data = 9'h090;
      591: data = 9'h08E;
      592: data = 9'h08C;
      593: data = 9'h08B;
      594: data = 9'h08A;
      595: data = 9'h089;
      596: data = 9'h088;
      597: data = 9'h088;
      598: data = 9'h088;
      599: data = 9'h089;
      600: data = 9'h089;
      601: data = 9'h089;
      602: data = 9'h08A;
      603: data = 9'h08B;
      604: data = 9'h08B;
      605: data = 9'h08C;
      606: data = 9'h08C;
      607: data = 9'h08C;
      608: data = 9'h08C;
      609: data = 9'h08B;
      610: data = 9'h08B;
      611: data = 9'h089;
      612: data = 9'h088;
      613: data = 9'h086;
      614: data = 9'h084;
      615: data = 9'h081;
      616: data = 9'h07E;
      617: data = 9'h07B;
      618: data = 9'h077;
      619: data = 9'h074;
      620: data = 9'h070;
      621: data = 9'h06C;
      622: data = 9'h069;
      623: data = 9'h065;
      624: data = 9'h062;
      625: data = 9'h05F;
      626: data = 9'h05C;
      627: data = 9'h05A;
      628: data = 9'h058;
      629: data = 9'h057;
      630: data = 9'h056;
      631: data = 9'h055;
      632: data = 9'h055;
      633: data = 9'h056;
      634: data = 9'h057;
      635: data = 9'h058;
      636: data = 9'h059;
      637: data = 9'h05B;
      638: data = 9'h05D;
      639: data = 9'h05F;
      640: data = 9'h061;
      641: data = 9'h063;
      642: data = 9'h064;
      643: data = 9'h065;
      644: data = 9'h066;
      645: data = 9'h066;
      646: data = 9'h066;
      647: data = 9'h064;
      648: data = 9'h063;
      649: data = 9'h060;
      650: data = 9'h05D;
      651: data = 9'h059;
      652: data = 9'h054;
      653: data = 9'h04F;
      654: data = 9'h049;
      655: data = 9'h043;
      656: data = 9'h03C;
      657: data = 9'h035;
      658: data = 9'h02F;
      659: data = 9'h028;
      660: data = 9'h022;
      661: data = 9'h01C;
      662: data = 9'h017;
      663: data = 9'h013;
      664: data = 9'h011;
      665: data = 9'h00F;
      666: data = 9'h00F;
      667: data = 9'h010;
      668: data = 9'h013;
      669: data = 9'h018;
      670: data = 9'h01F;
      671: data = 9'h028;
      672: data = 9'h032;
      673: data = 9'h03E;
      674: data = 9'h04D;
      675: data = 9'h05C;
      676: data = 9'h06E;
      677: data = 9'h081;
      678: data = 9'h095;
      679: data = 9'h0AA;
      680: data = 9'h0C1;
      681: data = 9'h0D8;
      682: data = 9'h0EF;
      683: data = 9'h106;
      684: data = 9'h11E;
      685: data = 9'h135;
      686: data = 9'h14B;
      687: data = 9'h161;
      688: data = 9'h175;
      689: data = 9'h189;
      690: data = 9'h19B;
      691: data = 9'h1AB;
      692: data = 9'h1BA;
      693: data = 9'h1C7;
      694: data = 9'h1D2;
      695: data = 9'h1DB;
      696: data = 9'h1E3;
      697: data = 9'h1E8;
      698: data = 9'h1EC;
      699: data = 9'h1EE;
      700: data = 9'h1EE;
      701: data = 9'h1ED;
      702: data = 9'h1EB;
      703: data = 9'h1E7;
      704: data = 9'h1E2;
      705: data = 9'h1DD;
      706: data = 9'h1D7;
      707: data = 9'h1D1;
      708: data = 9'h1CA;
      709: data = 9'h1C3;
      710: data = 9'h1BD;
      711: data = 9'h1B6;
      712: data = 9'h1B0;
      713: data = 9'h1AB;
      714: data = 9'h1A6;
      715: data = 9'h1A2;
      716: data = 9'h19E;
      717: data = 9'h19B;
      718: data = 9'h199;
      719: data = 9'h198;
      720: data = 9'h197;
      721: data = 9'h197;
      722: data = 9'h197;
      723: data = 9'h198;
      724: data = 9'h19A;
      725: data = 9'h19B;
      726: data = 9'h19D;
      727: data = 9'h19F;
      728: data = 9'h1A1;
      729: data = 9'h1A3;
      730: data = 9'h1A5;
      731: data = 9'h1A6;
      732: data = 9'h1A7;
      733: data = 9'h1A8;
      734: data = 9'h1A8;
      735: data = 9'h1A8;
      736: data = 9'h1A7;
      737: data = 9'h1A6;
      738: data = 9'h1A4;
      739: data = 9'h1A2;
      740: data = 9'h19F;
      741: data = 9'h19C;
      742: data = 9'h199;
      743: data = 9'h195;
      744: data = 9'h192;
      745: data = 9'h18E;
      746: data = 9'h18A;
      747: data = 9'h187;
      748: data = 9'h183;
      749: data = 9'h180;
      750: data = 9'h17D;
      751: data = 9'h17A;
      752: data = 9'h178;
      753: data = 9'h176;
      754: data = 9'h174;
      755: data = 9'h173;
      756: data = 9'h172;
      757: data = 9'h171;
      758: data = 9'h171;
      759: data = 9'h171;
      760: data = 9'h171;
      761: data = 9'h172;
      762: data = 9'h172;
      763: data = 9'h173;
      764: data = 9'h173;
      765: data = 9'h174;
      766: data = 9'h174;
      767: data = 9'h175;
      768: data = 9'h175;
      769: data = 9'h175;
      770: data = 9'h174;
      771: data = 9'h174;
      772: data = 9'h173;
      773: data = 9'h171;
      774: data = 9'h170;
      775: data = 9'h16E;
      776: data = 9'h16C;
      777: data = 9'h169;
      778: data = 9'h167;
      779: data = 9'h164;
      780: data = 9'h161;
      781: data = 9'h15E;
      782: data = 9'h15B;
      783: data = 9'h158;
      784: data = 9'h155;
      785: data = 9'h153;
      786: data = 9'h150;
      787: data = 9'h14E;
      788: data = 9'h14C;
      789: data = 9'h14A;
      790: data = 9'h148;
      791: data = 9'h147;
      792: data = 9'h146;
      793: data = 9'h145;
      794: data = 9'h145;
      795: data = 9'h144;
      796: data = 9'h144;
      797: data = 9'h144;
      798: data = 9'h144;
      799: data = 9'h144;
      800: data = 9'h145;
      801: data = 9'h145;
      802: data = 9'h145;
      803: data = 9'h145;
      804: data = 9'h145;
      805: data = 9'h144;
      806: data = 9'h144;
      807: data = 9'h143;
      808: data = 9'h142;
      809: data = 9'h140;
      810: data = 9'h13F;
      811: data = 9'h13D;
      812: data = 9'h13B;
      813: data = 9'h139;
      814: data = 9'h136;
      815: data = 9'h134;
      816: data = 9'h131;
      817: data = 9'h12F;
      818: data = 9'h12C;
      819: data = 9'h129;
      820: data = 9'h127;
      821: data = 9'h124;
      822: data = 9'h122;
      823: data = 9'h120;
      824: data = 9'h11E;
      825: data = 9'h11C;
      826: data = 9'h11A;
      827: data = 9'h119;
      828: data = 9'h118;
      829: data = 9'h117;
      830: data = 9'h117;
      831: data = 9'h116;
      832: data = 9'h116;
      833: data = 9'h116;
      834: data = 9'h116;
      835: data = 9'h116;
      836: data = 9'h116;
      837: data = 9'h116;
      838: data = 9'h116;
      839: data = 9'h116;
      840: data = 9'h115;
      841: data = 9'h115;
      842: data = 9'h114;
      843: data = 9'h113;
      844: data = 9'h112;
      845: data = 9'h111;
      846: data = 9'h10F;
      847: data = 9'h10D;
      848: data = 9'h10B;
      849: data = 9'h109;
      850: data = 9'h107;
      851: data = 9'h105;
      852: data = 9'h102;
      853: data = 9'h0FF;
      854: data = 9'h0FD;
      855: data = 9'h0FA;
      856: data = 9'h0F8;
      857: data = 9'h0F5;
      858: data = 9'h0F3;
      859: data = 9'h0F1;
      860: data = 9'h0EF;
      861: data = 9'h0ED;
      862: data = 9'h0EC;
      863: data = 9'h0EA;
      864: data = 9'h0E9;
      865: data = 9'h0E9;
      866: data = 9'h0E8;
      867: data = 9'h0E8;
      868: data = 9'h0E7;
      869: data = 9'h0E7;
      870: data = 9'h0E7;
      871: data = 9'h0E7;
      872: data = 9'h0E7;
      873: data = 9'h0E7;
      874: data = 9'h0E7;
      875: data = 9'h0E7;
      876: data = 9'h0E7;
      877: data = 9'h0E6;
      878: data = 9'h0E5;
      879: data = 9'h0E5;
      880: data = 9'h0E3;
      881: data = 9'h0E2;
      882: data = 9'h0E0;
      883: data = 9'h0DF;
      884: data = 9'h0DD;
      885: data = 9'h0DA;
      886: data = 9'h0D8;
      887: data = 9'h0D5;
      888: data = 9'h0D3;
      889: data = 9'h0D0;
      890: data = 9'h0CE;
      891: data = 9'h0CB;
      892: data = 9'h0C8;
      893: data = 9'h0C6;
      894: data = 9'h0C3;
      895: data = 9'h0C1;
      896: data = 9'h0BF;
      897: data = 9'h0BE;
      898: data = 9'h0BC;
      899: data = 9'h0BB;
      900: data = 9'h0BA;
      901: data = 9'h0B9;
      902: data = 9'h0B9;
      903: data = 9'h0B8;
      904: data = 9'h0B8;
      905: data = 9'h0B8;
      906: data = 9'h0B8;
      907: data = 9'h0B8;
      908: data = 9'h0B9;
      909: data = 9'h0B9;
      910: data = 9'h0B9;
      911: data = 9'h0B9;
      912: data = 9'h0B9;
      913: data = 9'h0B8;
      914: data = 9'h0B8;
      915: data = 9'h0B7;
      916: data = 9'h0B6;
      917: data = 9'h0B4;
      918: data = 9'h0B3;
      919: data = 9'h0B1;
      920: data = 9'h0AF;
      921: data = 9'h0AC;
      922: data = 9'h0AA;
      923: data = 9'h0A7;
      924: data = 9'h0A4;
      925: data = 9'h0A1;
      926: data = 9'h09E;
      927: data = 9'h09B;
      928: data = 9'h098;
      929: data = 9'h096;
      930: data = 9'h093;
      931: data = 9'h091;
      932: data = 9'h08F;
      933: data = 9'h08D;
      934: data = 9'h08B;
      935: data = 9'h08A;
      936: data = 9'h089;
      937: data = 9'h089;
      938: data = 9'h088;
      939: data = 9'h088;
      940: data = 9'h088;
      941: data = 9'h089;
      942: data = 9'h089;
      943: data = 9'h08A;
      944: data = 9'h08B;
      945: data = 9'h08B;
      946: data = 9'h08C;
      947: data = 9'h08C;
      948: data = 9'h08C;
      949: data = 9'h08C;
      950: data = 9'h08C;
      951: data = 9'h08B;
      952: data = 9'h08A;
      953: data = 9'h088;
      954: data = 9'h087;
      955: data = 9'h084;
      956: data = 9'h082;
      957: data = 9'h07F;
      958: data = 9'h07C;
      959: data = 9'h079;
      960: data = 9'h075;
      961: data = 9'h071;
      962: data = 9'h06E;
      963: data = 9'h06A;
      964: data = 9'h066;
      965: data = 9'h063;
      966: data = 9'h060;
      967: data = 9'h05D;
      968: data = 9'h05B;
      969: data = 9'h059;
      970: data = 9'h057;
      971: data = 9'h056;
      972: data = 9'h055;
      973: data = 9'h055;
      974: data = 9'h055;
      975: data = 9'h056;
      976: data = 9'h057;
      977: data = 9'h059;
      978: data = 9'h05B;
      979: data = 9'h05C;
      980: data = 9'h05E;
      981: data = 9'h060;
      982: data = 9'h062;
      983: data = 9'h064;
      984: data = 9'h065;
      985: data = 9'h066;
      986: data = 9'h066;
      987: data = 9'h066;
      988: data = 9'h065;
      989: data = 9'h063;
      990: data = 9'h061;
      991: data = 9'h05E;
      992: data = 9'h05A;
      993: data = 9'h056;
      994: data = 9'h051;
      995: data = 9'h04B;
      996: data = 9'h045;
      997: data = 9'h03E;
      998: data = 9'h038;
      999: data = 9'h031;
     1000: data = 9'h02A;
     1001: data = 9'h024;
     1002: data = 9'h01E;
     1003: data = 9'h019;
     1004: data = 9'h015;
     1005: data = 9'h011;
     1006: data = 9'h00F;
     1007: data = 9'h00F;
     1008: data = 9'h010;
     1009: data = 9'h012;
     1010: data = 9'h016;
     1011: data = 9'h01D;
     1012: data = 9'h025;
     1013: data = 9'h02E;
     1014: data = 9'h03A;
     1015: data = 9'h048;
     1016: data = 9'h057;
     1017: data = 9'h068;
     1018: data = 9'h07A;
     1019: data = 9'h08E;
     1020: data = 9'h0A3;
     1021: data = 9'h0B9;
     1022: data = 9'h0D0;
     1023: data = 9'h0E7;
    endcase
end

endmodule
