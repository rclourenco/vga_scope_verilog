module char_rom (
	input [10:0] address,
	output reg [7:0] data
);

always @(address)
begin
    case (address)
           0: data = 8'b00000000; //  0
           1: data = 8'b00000000; //  1
           2: data = 8'b00000000; //  2
           3: data = 8'b00000000; //  3
           4: data = 8'b00000000; //  4
           5: data = 8'b00000000; //  5
           6: data = 8'b00000000; //  6
           7: data = 8'b00000000; //  7
           8: data = 8'b00000000; //  8
           9: data = 8'b00000000; //  9
          10: data = 8'b00000000; //  a
          11: data = 8'b00000000; //  b
          12: data = 8'b00000000; //  c
          13: data = 8'b00000000; //  d
          14: data = 8'b00000000; //  e
          15: data = 8'b00000000; //  f
          //    code x01
          16: data = 8'b00000000; //  0
          17: data = 8'b00000000; //  1
          18: data = 8'b01111110; //  2  ******
          19: data = 8'b10000001; //  3 *      *
          20: data = 8'b10100101; //  4 * *  * *
          21: data = 8'b10000001; //  5 *      *
          22: data = 8'b10000001; //  6 *      *
          23: data = 8'b10111101; //  7 * **** *
          24: data = 8'b10011001; //  8 *  **  *
          25: data = 8'b10000001; //  9 *      *
          26: data = 8'b10000001; //  a *      *
          27: data = 8'b01111110; //  b  ******
          28: data = 8'b00000000; //  c
          29: data = 8'b00000000; //  d
          30: data = 8'b00000000; //  e
          31: data = 8'b00000000; //  f
          //    code x02
          32: data = 8'b00000000; //  0
          33: data = 8'b00000000; //  1
          34: data = 8'b01111110; //  2  ******
          35: data = 8'b11111111; //  3 ********
          36: data = 8'b11011011; //  4 ** ** **
          37: data = 8'b11111111; //  5 ********
          38: data = 8'b11111111; //  6 ********
          39: data = 8'b11000011; //  7 **    **
          40: data = 8'b11100111; //  8 ***  ***
          41: data = 8'b11111111; //  9 ********
          42: data = 8'b11111111; //  a ********
          43: data = 8'b01111110; //  b  ******
          44: data = 8'b00000000; //  c
          45: data = 8'b00000000; //  d
          46: data = 8'b00000000; //  e
          47: data = 8'b00000000; //  f
          //    code x03
          48: data = 8'b00000000; //  0
          49: data = 8'b00000000; //  1
          50: data = 8'b00000000; //  2
          51: data = 8'b00000000; //  3
          52: data = 8'b01101100; //  4  ** **
          53: data = 8'b11111110; //  5 *******
          54: data = 8'b11111110; //  6 *******
          55: data = 8'b11111110; //  7 *******
          56: data = 8'b11111110; //  8 *******
          57: data = 8'b01111100; //  9  *****
          58: data = 8'b00111000; //  a   ***
          59: data = 8'b00010000; //  b    *
          60: data = 8'b00000000; //  c
          61: data = 8'b00000000; //  d
          62: data = 8'b00000000; //  e
          63: data = 8'b00000000; //  f
          //    code x04
          64: data = 8'b00000000; //  0
          65: data = 8'b00000000; //  1
          66: data = 8'b00000000; //  2
          67: data = 8'b00000000; //  3
          68: data = 8'b00010000; //  4    *
          69: data = 8'b00111000; //  5   ***
          70: data = 8'b01111100; //  6  *****
          71: data = 8'b11111110; //  7 *******
          72: data = 8'b01111100; //  8  *****
          73: data = 8'b00111000; //  9   ***
          74: data = 8'b00010000; //  a    *
          75: data = 8'b00000000; //  b
          76: data = 8'b00000000; //  c
          77: data = 8'b00000000; //  d
          78: data = 8'b00000000; //  e
          79: data = 8'b00000000; //  f
          //    code x05
          80: data = 8'b00000000; //  0
          81: data = 8'b00000000; //  1
          82: data = 8'b00000000; //  2
          83: data = 8'b00011000; //  3    **
          84: data = 8'b00111100; //  4   ****
          85: data = 8'b00111100; //  5   ****
          86: data = 8'b11100111; //  6 ***  ***
          87: data = 8'b11100111; //  7 ***  ***
          88: data = 8'b11100111; //  8 ***  ***
          89: data = 8'b00011000; //  9    **
          90: data = 8'b00011000; //  a    **
          91: data = 8'b00111100; //  b   ****
          92: data = 8'b00000000; //  c
          93: data = 8'b00000000; //  d
          94: data = 8'b00000000; //  e
          95: data = 8'b00000000; //  f
          //    code x06
          96: data = 8'b00000000; //  0
          97: data = 8'b00000000; //  1
          98: data = 8'b00000000; //  2
          99: data = 8'b00011000; //  3    **
         100: data = 8'b00111100; //  4   ****
         101: data = 8'b01111110; //  5  ******
         102: data = 8'b11111111; //  6 ********
         103: data = 8'b11111111; //  7 ********
         104: data = 8'b01111110; //  8  ******
         105: data = 8'b00011000; //  9    **
         106: data = 8'b00011000; //  a    **
         107: data = 8'b00111100; //  b   ****
         108: data = 8'b00000000; //  c
         109: data = 8'b00000000; //  d
         110: data = 8'b00000000; //  e
         111: data = 8'b00000000; //  f
          //    code x07
         112: data = 8'b00000000; //  0
         113: data = 8'b00000000; //  1
         114: data = 8'b00000000; //  2
         115: data = 8'b00000000; //  3
         116: data = 8'b00000000; //  4
         117: data = 8'b00000000; //  5
         118: data = 8'b00011000; //  6    **
         119: data = 8'b00111100; //  7   ****
         120: data = 8'b00111100; //  8   ****
         121: data = 8'b00011000; //  9    **
         122: data = 8'b00000000; //  a
         123: data = 8'b00000000; //  b
         124: data = 8'b00000000; //  c
         125: data = 8'b00000000; //  d
         126: data = 8'b00000000; //  e
         127: data = 8'b00000000; //  f
          //    code x08
         128: data = 8'b11111111; //  0 ********
         129: data = 8'b11111111; //  1 ********
         130: data = 8'b11111111; //  2 ********
         131: data = 8'b11111111; //  3 ********
         132: data = 8'b11111111; //  4 ********
         133: data = 8'b11111111; //  5 ********
         134: data = 8'b11100111; //  6 ***  ***
         135: data = 8'b11000011; //  7 **    **
         136: data = 8'b11000011; //  8 **    **
         137: data = 8'b11100111; //  9 ***  ***
         138: data = 8'b11111111; //  a ********
         139: data = 8'b11111111; //  b ********
         140: data = 8'b11111111; //  c ********
         141: data = 8'b11111111; //  d ********
         142: data = 8'b11111111; //  e ********
         143: data = 8'b11111111; //  f ********
          //    code x09
         144: data = 8'b00000000; //  0
         145: data = 8'b00000000; //  1
         146: data = 8'b00000000; //  2
         147: data = 8'b00000000; //  3
         148: data = 8'b00000000; //  4
         149: data = 8'b00111100; //  5   ****
         150: data = 8'b01100110; //  6  **  **
         151: data = 8'b01000010; //  7  *    *
         152: data = 8'b01000010; //  8  *    *
         153: data = 8'b01100110; //  9  **  **
         154: data = 8'b00111100; //  a   ****
         155: data = 8'b00000000; //  b
         156: data = 8'b00000000; //  c
         157: data = 8'b00000000; //  d
         158: data = 8'b00000000; //  e
         159: data = 8'b00000000; //  f
          //    code x0a
         160: data = 8'b11111111; //  0 ********
         161: data = 8'b11111111; //  1 ********
         162: data = 8'b11111111; //  2 ********
         163: data = 8'b11111111; //  3 ********
         164: data = 8'b11111111; //  4 ********
         165: data = 8'b11000011; //  5 **    **
         166: data = 8'b10011001; //  6 *  **  *
         167: data = 8'b10111101; //  7 * **** *
         168: data = 8'b10111101; //  8 * **** *
         169: data = 8'b10011001; //  9 *  **  *
         170: data = 8'b11000011; //  a **    **
         171: data = 8'b11111111; //  b ********
         172: data = 8'b11111111; //  c ********
         173: data = 8'b11111111; //  d ********
         174: data = 8'b11111111; //  e ********
         175: data = 8'b11111111; //  f ********
          //    code x0b
         176: data = 8'b00000000; //  0
         177: data = 8'b00000000; //  1
         178: data = 8'b00011110; //  2    ****
         179: data = 8'b00001110; //  3     ***
         180: data = 8'b00011010; //  4    ** *
         181: data = 8'b00110010; //  5   **  *
         182: data = 8'b01111000; //  6  ****
         183: data = 8'b11001100; //  7 **  **
         184: data = 8'b11001100; //  8 **  **
         185: data = 8'b11001100; //  9 **  **
         186: data = 8'b11001100; //  a **  **
         187: data = 8'b01111000; //  b  ****
         188: data = 8'b00000000; //  c
         189: data = 8'b00000000; //  d
         190: data = 8'b00000000; //  e
         191: data = 8'b00000000; //  f
          //    code x0c
         192: data = 8'b00000000; //  0
         193: data = 8'b00000000; //  1
         194: data = 8'b00111100; //  2   ****
         195: data = 8'b01100110; //  3  **  **
         196: data = 8'b01100110; //  4  **  **
         197: data = 8'b01100110; //  5  **  **
         198: data = 8'b01100110; //  6  **  **
         199: data = 8'b00111100; //  7   ****
         200: data = 8'b00011000; //  8    **
         201: data = 8'b01111110; //  9  ******
         202: data = 8'b00011000; //  a    **
         203: data = 8'b00011000; //  b    **
         204: data = 8'b00000000; //  c
         205: data = 8'b00000000; //  d
         206: data = 8'b00000000; //  e
         207: data = 8'b00000000; //  f
          //    code x0d
         208: data = 8'b00000000; //  0
         209: data = 8'b00000000; //  1
         210: data = 8'b00111111; //  2   ******
         211: data = 8'b00110011; //  3   **  **
         212: data = 8'b00111111; //  4   ******
         213: data = 8'b00110000; //  5   **
         214: data = 8'b00110000; //  6   **
         215: data = 8'b00110000; //  7   **
         216: data = 8'b00110000; //  8   **
         217: data = 8'b01110000; //  9  ***
         218: data = 8'b11110000; //  a ****
         219: data = 8'b11100000; //  b ***
         220: data = 8'b00000000; //  c
         221: data = 8'b00000000; //  d
         222: data = 8'b00000000; //  e
         223: data = 8'b00000000; //  f
          //    code x0e
         224: data = 8'b00000000; //  0
         225: data = 8'b00000000; //  1
         226: data = 8'b01111111; //  2  *******
         227: data = 8'b01100011; //  3  **   **
         228: data = 8'b01111111; //  4  *******
         229: data = 8'b01100011; //  5  **   **
         230: data = 8'b01100011; //  6  **   **
         231: data = 8'b01100011; //  7  **   **
         232: data = 8'b01100011; //  8  **   **
         233: data = 8'b01100111; //  9  **  ***
         234: data = 8'b11100111; //  a ***  ***
         235: data = 8'b11100110; //  b ***  **
         236: data = 8'b11000000; //  c **
         237: data = 8'b00000000; //  d
         238: data = 8'b00000000; //  e
         239: data = 8'b00000000; //  f
          //    code x0f
         240: data = 8'b00000000; //  0
         241: data = 8'b00000000; //  1
         242: data = 8'b00000000; //  2
         243: data = 8'b00011000; //  3    **
         244: data = 8'b00011000; //  4    **
         245: data = 8'b11011011; //  5 ** ** **
         246: data = 8'b00111100; //  6   ****
         247: data = 8'b11100111; //  7 ***  ***
         248: data = 8'b00111100; //  8   ****
         249: data = 8'b11011011; //  9 ** ** **
         250: data = 8'b00011000; //  a    **
         251: data = 8'b00011000; //  b    **
         252: data = 8'b00000000; //  c
         253: data = 8'b00000000; //  d
         254: data = 8'b00000000; //  e
         255: data = 8'b00000000; //  f
          //    code x10
         256: data = 8'b00000000; //  0
         257: data = 8'b10000000; //  1 *
         258: data = 8'b11000000; //  2 **
         259: data = 8'b11100000; //  3 ***
         260: data = 8'b11110000; //  4 ****
         261: data = 8'b11111000; //  5 *****
         262: data = 8'b11111110; //  6 *******
         263: data = 8'b11111000; //  7 *****
         264: data = 8'b11110000; //  8 ****
         265: data = 8'b11100000; //  9 ***
         266: data = 8'b11000000; //  a **
         267: data = 8'b10000000; //  b *
         268: data = 8'b00000000; //  c
         269: data = 8'b00000000; //  d
         270: data = 8'b00000000; //  e
         271: data = 8'b00000000; //  f
          //    code x11
         272: data = 8'b00000000; //  0
         273: data = 8'b00000010; //  1       *
         274: data = 8'b00000110; //  2      **
         275: data = 8'b00001110; //  3     ***
         276: data = 8'b00011110; //  4    ****
         277: data = 8'b00111110; //  5   *****
         278: data = 8'b11111110; //  6 *******
         279: data = 8'b00111110; //  7   *****
         280: data = 8'b00011110; //  8    ****
         281: data = 8'b00001110; //  9     ***
         282: data = 8'b00000110; //  a      **
         283: data = 8'b00000010; //  b       *
         284: data = 8'b00000000; //  c
         285: data = 8'b00000000; //  d
         286: data = 8'b00000000; //  e
         287: data = 8'b00000000; //  f
          //    code x12
         288: data = 8'b00000000; //  0
         289: data = 8'b00000000; //  1
         290: data = 8'b00011000; //  2    **
         291: data = 8'b00111100; //  3   ****
         292: data = 8'b01111110; //  4  ******
         293: data = 8'b00011000; //  5    **
         294: data = 8'b00011000; //  6    **
         295: data = 8'b00011000; //  7    **
         296: data = 8'b01111110; //  8  ******
         297: data = 8'b00111100; //  9   ****
         298: data = 8'b00011000; //  a    **
         299: data = 8'b00000000; //  b
         300: data = 8'b00000000; //  c
         301: data = 8'b00000000; //  d
         302: data = 8'b00000000; //  e
         303: data = 8'b00000000; //  f
          //    code x13
         304: data = 8'b00000000; //  0
         305: data = 8'b00000000; //  1
         306: data = 8'b01100110; //  2  **  **
         307: data = 8'b01100110; //  3  **  **
         308: data = 8'b01100110; //  4  **  **
         309: data = 8'b01100110; //  5  **  **
         310: data = 8'b01100110; //  6  **  **
         311: data = 8'b01100110; //  7  **  **
         312: data = 8'b01100110; //  8  **  **
         313: data = 8'b00000000; //  9
         314: data = 8'b01100110; //  a  **  **
         315: data = 8'b01100110; //  b  **  **
         316: data = 8'b00000000; //  c
         317: data = 8'b00000000; //  d
         318: data = 8'b00000000; //  e
         319: data = 8'b00000000; //  f
          //    code x14
         320: data = 8'b00000000; //  0
         321: data = 8'b00000000; //  1
         322: data = 8'b01111111; //  2  *******
         323: data = 8'b11011011; //  3 ** ** **
         324: data = 8'b11011011; //  4 ** ** **
         325: data = 8'b11011011; //  5 ** ** **
         326: data = 8'b01111011; //  6  **** **
         327: data = 8'b00011011; //  7    ** **
         328: data = 8'b00011011; //  8    ** **
         329: data = 8'b00011011; //  9    ** **
         330: data = 8'b00011011; //  a    ** **
         331: data = 8'b00011011; //  b    ** **
         332: data = 8'b00000000; //  c
         333: data = 8'b00000000; //  d
         334: data = 8'b00000000; //  e
         335: data = 8'b00000000; //  f
          //    code x15
         336: data = 8'b00000000; //  0
         337: data = 8'b01111100; //  1  *****
         338: data = 8'b11000110; //  2 **   **
         339: data = 8'b01100000; //  3  **
         340: data = 8'b00111000; //  4   ***
         341: data = 8'b01101100; //  5  ** **
         342: data = 8'b11000110; //  6 **   **
         343: data = 8'b11000110; //  7 **   **
         344: data = 8'b01101100; //  8  ** **
         345: data = 8'b00111000; //  9   ***
         346: data = 8'b00001100; //  a     **
         347: data = 8'b11000110; //  b **   **
         348: data = 8'b01111100; //  c  *****
         349: data = 8'b00000000; //  d
         350: data = 8'b00000000; //  e
         351: data = 8'b00000000; //  f
          //    code x16
         352: data = 8'b00000000; //  0
         353: data = 8'b00000000; //  1
         354: data = 8'b00000000; //  2
         355: data = 8'b00000000; //  3
         356: data = 8'b00000000; //  4
         357: data = 8'b00000000; //  5
         358: data = 8'b00000000; //  6
         359: data = 8'b00000000; //  7
         360: data = 8'b11111110; //  8 *******
         361: data = 8'b11111110; //  9 *******
         362: data = 8'b11111110; //  a *******
         363: data = 8'b11111110; //  b *******
         364: data = 8'b00000000; //  c
         365: data = 8'b00000000; //  d
         366: data = 8'b00000000; //  e
         367: data = 8'b00000000; //  f
          //    code x17
         368: data = 8'b00000000; //  0
         369: data = 8'b00000000; //  1
         370: data = 8'b00011000; //  2    **
         371: data = 8'b00111100; //  3   ****
         372: data = 8'b01111110; //  4  ******
         373: data = 8'b00011000; //  5    **
         374: data = 8'b00011000; //  6    **
         375: data = 8'b00011000; //  7    **
         376: data = 8'b01111110; //  8  ******
         377: data = 8'b00111100; //  9   ****
         378: data = 8'b00011000; //  a    **
         379: data = 8'b01111110; //  b  ******
         380: data = 8'b00110000; //  c
         381: data = 8'b00000000; //  d
         382: data = 8'b00000000; //  e
         383: data = 8'b00000000; //  f
          //    code x18
         384: data = 8'b00000000; //  0
         385: data = 8'b00000000; //  1
         386: data = 8'b00011000; //  2    **
         387: data = 8'b00111100; //  3   ****
         388: data = 8'b01111110; //  4  ******
         389: data = 8'b00011000; //  5    **
         390: data = 8'b00011000; //  6    **
         391: data = 8'b00011000; //  7    **
         392: data = 8'b00011000; //  8    **
         393: data = 8'b00011000; //  9    **
         394: data = 8'b00011000; //  a    **
         395: data = 8'b00011000; //  b    **
         396: data = 8'b00000000; //  c
         397: data = 8'b00000000; //  d
         398: data = 8'b00000000; //  e
         399: data = 8'b00000000; //  f
          //    code x19
         400: data = 8'b00000000; //  0
         401: data = 8'b00000000; //  1
         402: data = 8'b00011000; //  2    **
         403: data = 8'b00011000; //  3    **
         404: data = 8'b00011000; //  4    **
         405: data = 8'b00011000; //  5    **
         406: data = 8'b00011000; //  6    **
         407: data = 8'b00011000; //  7    **
         408: data = 8'b00011000; //  8    **
         409: data = 8'b01111110; //  9  ******
         410: data = 8'b00111100; //  a   ****
         411: data = 8'b00011000; //  b    **
         412: data = 8'b00000000; //  c
         413: data = 8'b00000000; //  d
         414: data = 8'b00000000; //  e
         415: data = 8'b00000000; //  f
          //    code x1a
         416: data = 8'b00000000; //  0
         417: data = 8'b00000000; //  1
         418: data = 8'b00000000; //  2
         419: data = 8'b00000000; //  3
         420: data = 8'b00000000; //  4
         421: data = 8'b00011000; //  5    **
         422: data = 8'b00001100; //  6     **
         423: data = 8'b11111110; //  7 *******
         424: data = 8'b00001100; //  8     **
         425: data = 8'b00011000; //  9    **
         426: data = 8'b00000000; //  a
         427: data = 8'b00000000; //  b
         428: data = 8'b00000000; //  c
         429: data = 8'b00000000; //  d
         430: data = 8'b00000000; //  e
         431: data = 8'b00000000; //  f
          //    code x1b
         432: data = 8'b00000000; //  0
         433: data = 8'b00000000; //  1
         434: data = 8'b00000000; //  2
         435: data = 8'b00000000; //  3
         436: data = 8'b00000000; //  4
         437: data = 8'b00110000; //  5   **
         438: data = 8'b01100000; //  6  **
         439: data = 8'b11111110; //  7 *******
         440: data = 8'b01100000; //  8  **
         441: data = 8'b00110000; //  9   **
         442: data = 8'b00000000; //  a
         443: data = 8'b00000000; //  b
         444: data = 8'b00000000; //  c
         445: data = 8'b00000000; //  d
         446: data = 8'b00000000; //  e
         447: data = 8'b00000000; //  f
          //    code x1c
         448: data = 8'b00000000; //  0
         449: data = 8'b00000000; //  1
         450: data = 8'b00000000; //  2
         451: data = 8'b00000000; //  3
         452: data = 8'b00000000; //  4
         453: data = 8'b00000000; //  5
         454: data = 8'b11000000; //  6 **
         455: data = 8'b11000000; //  7 **
         456: data = 8'b11000000; //  8 **
         457: data = 8'b11111110; //  9 *******
         458: data = 8'b00000000; //  a
         459: data = 8'b00000000; //  b
         460: data = 8'b00000000; //  c
         461: data = 8'b00000000; //  d
         462: data = 8'b00000000; //  e
         463: data = 8'b00000000; //  f
          //    code x1d
         464: data = 8'b00000000; //  0
         465: data = 8'b00000000; //  1
         466: data = 8'b00000000; //  2
         467: data = 8'b00000000; //  3
         468: data = 8'b00000000; //  4
         469: data = 8'b00100100; //  5   *  *
         470: data = 8'b01100110; //  6  **  **
         471: data = 8'b11111111; //  7 ********
         472: data = 8'b01100110; //  8  **  **
         473: data = 8'b00100100; //  9   *  *
         474: data = 8'b00000000; //  a
         475: data = 8'b00000000; //  b
         476: data = 8'b00000000; //  c
         477: data = 8'b00000000; //  d
         478: data = 8'b00000000; //  e
         479: data = 8'b00000000; //  f
          //    code x1e
         480: data = 8'b00000000; //  0
         481: data = 8'b00000000; //  1
         482: data = 8'b00000000; //  2
         483: data = 8'b00000000; //  3
         484: data = 8'b00010000; //  4    *
         485: data = 8'b00111000; //  5   ***
         486: data = 8'b00111000; //  6   ***
         487: data = 8'b01111100; //  7  *****
         488: data = 8'b01111100; //  8  *****
         489: data = 8'b11111110; //  9 *******
         490: data = 8'b11111110; //  a *******
         491: data = 8'b00000000; //  b
         492: data = 8'b00000000; //  c
         493: data = 8'b00000000; //  d
         494: data = 8'b00000000; //  e
         495: data = 8'b00000000; //  f
          //    code x1f
         496: data = 8'b00000000; //  0
         497: data = 8'b00000000; //  1
         498: data = 8'b00000000; //  2
         499: data = 8'b00000000; //  3
         500: data = 8'b11111110; //  4 *******
         501: data = 8'b11111110; //  5 *******
         502: data = 8'b01111100; //  6  *****
         503: data = 8'b01111100; //  7  *****
         504: data = 8'b00111000; //  8   ***
         505: data = 8'b00111000; //  9   ***
         506: data = 8'b00010000; //  a    *
         507: data = 8'b00000000; //  b
         508: data = 8'b00000000; //  c
         509: data = 8'b00000000; //  d
         510: data = 8'b00000000; //  e
         511: data = 8'b00000000; //  f
          //    code x20
         512: data = 8'b00000000; //  0
         513: data = 8'b00000000; //  1
         514: data = 8'b00000000; //  2
         515: data = 8'b00000000; //  3
         516: data = 8'b00000000; //  4
         517: data = 8'b00000000; //  5
         518: data = 8'b00000000; //  6
         519: data = 8'b00000000; //  7
         520: data = 8'b00000000; //  8
         521: data = 8'b00000000; //  9
         522: data = 8'b00000000; //  a
         523: data = 8'b00000000; //  b
         524: data = 8'b00000000; //  c
         525: data = 8'b00000000; //  d
         526: data = 8'b00000000; //  e
         527: data = 8'b00000000; //  f
          //    code x21
         528: data = 8'b00000000; //  0
         529: data = 8'b00000000; //  1
         530: data = 8'b00011000; //  2    **
         531: data = 8'b00111100; //  3   ****
         532: data = 8'b00111100; //  4   ****
         533: data = 8'b00111100; //  5   ****
         534: data = 8'b00011000; //  6    **
         535: data = 8'b00011000; //  7    **
         536: data = 8'b00011000; //  8    **
         537: data = 8'b00000000; //  9
         538: data = 8'b00011000; //  a    **
         539: data = 8'b00011000; //  b    **
         540: data = 8'b00000000; //  c
         541: data = 8'b00000000; //  d
         542: data = 8'b00000000; //  e
         543: data = 8'b00000000; //  f
          //    code x22
         544: data = 8'b00000000; //  0
         545: data = 8'b01100110; //  1  **  **
         546: data = 8'b01100110; //  2  **  **
         547: data = 8'b01100110; //  3  **  **
         548: data = 8'b00100100; //  4   *  *
         549: data = 8'b00000000; //  5
         550: data = 8'b00000000; //  6
         551: data = 8'b00000000; //  7
         552: data = 8'b00000000; //  8
         553: data = 8'b00000000; //  9
         554: data = 8'b00000000; //  a
         555: data = 8'b00000000; //  b
         556: data = 8'b00000000; //  c
         557: data = 8'b00000000; //  d
         558: data = 8'b00000000; //  e
         559: data = 8'b00000000; //  f
          //    code x23
         560: data = 8'b00000000; //  0
         561: data = 8'b00000000; //  1
         562: data = 8'b00000000; //  2
         563: data = 8'b01101100; //  3  ** **
         564: data = 8'b01101100; //  4  ** **
         565: data = 8'b11111110; //  5 *******
         566: data = 8'b01101100; //  6  ** **
         567: data = 8'b01101100; //  7  ** **
         568: data = 8'b01101100; //  8  ** **
         569: data = 8'b11111110; //  9 *******
         570: data = 8'b01101100; //  a  ** **
         571: data = 8'b01101100; //  b  ** **
         572: data = 8'b00000000; //  c
         573: data = 8'b00000000; //  d
         574: data = 8'b00000000; //  e
         575: data = 8'b00000000; //  f
          //    code x24
         576: data = 8'b00011000; //  0     **
         577: data = 8'b00011000; //  1     **
         578: data = 8'b01111100; //  2   *****
         579: data = 8'b11000110; //  3  **   **
         580: data = 8'b11000010; //  4  **    *
         581: data = 8'b11000000; //  5  **
         582: data = 8'b01111100; //  6   *****
         583: data = 8'b00000110; //  7       **
         584: data = 8'b00000110; //  8       **
         585: data = 8'b10000110; //  9  *    **
         586: data = 8'b11000110; //  a  **   **
         587: data = 8'b01111100; //  b   *****
         588: data = 8'b00011000; //  c     **
         589: data = 8'b00011000; //  d     **
         590: data = 8'b00000000; //  e
         591: data = 8'b00000000; //  f
          //    code x25
         592: data = 8'b00000000; //  0
         593: data = 8'b00000000; //  1
         594: data = 8'b00000000; //  2
         595: data = 8'b00000000; //  3
         596: data = 8'b11000010; //  4 **    *
         597: data = 8'b11000110; //  5 **   **
         598: data = 8'b00001100; //  6     **
         599: data = 8'b00011000; //  7    **
         600: data = 8'b00110000; //  8   **
         601: data = 8'b01100000; //  9  **
         602: data = 8'b11000110; //  a **   **
         603: data = 8'b10000110; //  b *    **
         604: data = 8'b00000000; //  c
         605: data = 8'b00000000; //  d
         606: data = 8'b00000000; //  e
         607: data = 8'b00000000; //  f
          //    code x26
         608: data = 8'b00000000; //  0
         609: data = 8'b00000000; //  1
         610: data = 8'b00111000; //  2   ***
         611: data = 8'b01101100; //  3  ** **
         612: data = 8'b01101100; //  4  ** **
         613: data = 8'b00111000; //  5   ***
         614: data = 8'b01110110; //  6  *** **
         615: data = 8'b11011100; //  7 ** ***
         616: data = 8'b11001100; //  8 **  **
         617: data = 8'b11001100; //  9 **  **
         618: data = 8'b11001100; //  a **  **
         619: data = 8'b01110110; //  b  *** **
         620: data = 8'b00000000; //  c
         621: data = 8'b00000000; //  d
         622: data = 8'b00000000; //  e
         623: data = 8'b00000000; //  f
          //    code x27
         624: data = 8'b00000000; //  0
         625: data = 8'b00110000; //  1   **
         626: data = 8'b00110000; //  2   **
         627: data = 8'b00110000; //  3   **
         628: data = 8'b01100000; //  4  **
         629: data = 8'b00000000; //  5
         630: data = 8'b00000000; //  6
         631: data = 8'b00000000; //  7
         632: data = 8'b00000000; //  8
         633: data = 8'b00000000; //  9
         634: data = 8'b00000000; //  a
         635: data = 8'b00000000; //  b
         636: data = 8'b00000000; //  c
         637: data = 8'b00000000; //  d
         638: data = 8'b00000000; //  e
         639: data = 8'b00000000; //  f
          //    code x28
         640: data = 8'b00000000; //  0
         641: data = 8'b00000000; //  1
         642: data = 8'b00001100; //  2     **
         643: data = 8'b00011000; //  3    **
         644: data = 8'b00110000; //  4   **
         645: data = 8'b00110000; //  5   **
         646: data = 8'b00110000; //  6   **
         647: data = 8'b00110000; //  7   **
         648: data = 8'b00110000; //  8   **
         649: data = 8'b00110000; //  9   **
         650: data = 8'b00011000; //  a    **
         651: data = 8'b00001100; //  b     **
         652: data = 8'b00000000; //  c
         653: data = 8'b00000000; //  d
         654: data = 8'b00000000; //  e
         655: data = 8'b00000000; //  f
          //    code x29
         656: data = 8'b00000000; //  0
         657: data = 8'b00000000; //  1
         658: data = 8'b00110000; //  2   **
         659: data = 8'b00011000; //  3    **
         660: data = 8'b00001100; //  4     **
         661: data = 8'b00001100; //  5     **
         662: data = 8'b00001100; //  6     **
         663: data = 8'b00001100; //  7     **
         664: data = 8'b00001100; //  8     **
         665: data = 8'b00001100; //  9     **
         666: data = 8'b00011000; //  a    **
         667: data = 8'b00110000; //  b   **
         668: data = 8'b00000000; //  c
         669: data = 8'b00000000; //  d
         670: data = 8'b00000000; //  e
         671: data = 8'b00000000; //  f
          //    code x2a
         672: data = 8'b00000000; //  0
         673: data = 8'b00000000; //  1
         674: data = 8'b00000000; //  2
         675: data = 8'b00000000; //  3
         676: data = 8'b00000000; //  4
         677: data = 8'b01100110; //  5  **  **
         678: data = 8'b00111100; //  6   ****
         679: data = 8'b11111111; //  7 ********
         680: data = 8'b00111100; //  8   ****
         681: data = 8'b01100110; //  9  **  **
         682: data = 8'b00000000; //  a
         683: data = 8'b00000000; //  b
         684: data = 8'b00000000; //  c
         685: data = 8'b00000000; //  d
         686: data = 8'b00000000; //  e
         687: data = 8'b00000000; //  f
          //    code x2b
         688: data = 8'b00000000; //  0
         689: data = 8'b00000000; //  1
         690: data = 8'b00000000; //  2
         691: data = 8'b00000000; //  3
         692: data = 8'b00000000; //  4
         693: data = 8'b00011000; //  5    **
         694: data = 8'b00011000; //  6    **
         695: data = 8'b01111110; //  7  ******
         696: data = 8'b00011000; //  8    **
         697: data = 8'b00011000; //  9    **
         698: data = 8'b00000000; //  a
         699: data = 8'b00000000; //  b
         700: data = 8'b00000000; //  c
         701: data = 8'b00000000; //  d
         702: data = 8'b00000000; //  e
         703: data = 8'b00000000; //  f
          //    code x2c
         704: data = 8'b00000000; //  0
         705: data = 8'b00000000; //  1
         706: data = 8'b00000000; //  2
         707: data = 8'b00000000; //  3
         708: data = 8'b00000000; //  4
         709: data = 8'b00000000; //  5
         710: data = 8'b00000000; //  6
         711: data = 8'b00000000; //  7
         712: data = 8'b00000000; //  8
         713: data = 8'b00011000; //  9    **
         714: data = 8'b00011000; //  a    **
         715: data = 8'b00011000; //  b    **
         716: data = 8'b00110000; //  c   **
         717: data = 8'b00000000; //  d
         718: data = 8'b00000000; //  e
         719: data = 8'b00000000; //  f
          //    code x2d
         720: data = 8'b00000000; //  0
         721: data = 8'b00000000; //  1
         722: data = 8'b00000000; //  2
         723: data = 8'b00000000; //  3
         724: data = 8'b00000000; //  4
         725: data = 8'b00000000; //  5
         726: data = 8'b00000000; //  6
         727: data = 8'b01111110; //  7  ******
         728: data = 8'b00000000; //  8
         729: data = 8'b00000000; //  9
         730: data = 8'b00000000; //  a
         731: data = 8'b00000000; //  b
         732: data = 8'b00000000; //  c
         733: data = 8'b00000000; //  d
         734: data = 8'b00000000; //  e
         735: data = 8'b00000000; //  f
          //    code x2e
         736: data = 8'b00000000; //  0
         737: data = 8'b00000000; //  1
         738: data = 8'b00000000; //  2
         739: data = 8'b00000000; //  3
         740: data = 8'b00000000; //  4
         741: data = 8'b00000000; //  5
         742: data = 8'b00000000; //  6
         743: data = 8'b00000000; //  7
         744: data = 8'b00000000; //  8
         745: data = 8'b00000000; //  9
         746: data = 8'b00011000; //  a    **
         747: data = 8'b00011000; //  b    **
         748: data = 8'b00000000; //  c
         749: data = 8'b00000000; //  d
         750: data = 8'b00000000; //  e
         751: data = 8'b00000000; //  f
          //    code x2f
         752: data = 8'b00000000; //  0
         753: data = 8'b00000000; //  1
         754: data = 8'b00000000; //  2
         755: data = 8'b00000000; //  3
         756: data = 8'b00000010; //  4       *
         757: data = 8'b00000110; //  5      **
         758: data = 8'b00001100; //  6     **
         759: data = 8'b00011000; //  7    **
         760: data = 8'b00110000; //  8   **
         761: data = 8'b01100000; //  9  **
         762: data = 8'b11000000; //  a **
         763: data = 8'b10000000; //  b *
         764: data = 8'b00000000; //  c
         765: data = 8'b00000000; //  d
         766: data = 8'b00000000; //  e
         767: data = 8'b00000000; //  f
          //    code x30
         768: data = 8'b00000000; //  0
         769: data = 8'b00000000; //  1
         770: data = 8'b01111100; //  2  *****
         771: data = 8'b11000110; //  3 **   **
         772: data = 8'b11000110; //  4 **   **
         773: data = 8'b11001110; //  5 **  ***
         774: data = 8'b11011110; //  6 ** ****
         775: data = 8'b11110110; //  7 **** **
         776: data = 8'b11100110; //  8 ***  **
         777: data = 8'b11000110; //  9 **   **
         778: data = 8'b11000110; //  a **   **
         779: data = 8'b01111100; //  b  *****
         780: data = 8'b00000000; //  c
         781: data = 8'b00000000; //  d
         782: data = 8'b00000000; //  e
         783: data = 8'b00000000; //  f
          //    code x31
         784: data = 8'b00000000; //  0
         785: data = 8'b00000000; //  1
         786: data = 8'b00011000; //  2
         787: data = 8'b00111000; //  3
         788: data = 8'b01111000; //  4    **
         789: data = 8'b00011000; //  5   ***
         790: data = 8'b00011000; //  6  ****
         791: data = 8'b00011000; //  7    **
         792: data = 8'b00011000; //  8    **
         793: data = 8'b00011000; //  9    **
         794: data = 8'b00011000; //  a    **
         795: data = 8'b01111110; //  b    **
         796: data = 8'b00000000; //  c    **
         797: data = 8'b00000000; //  d  ******
         798: data = 8'b00000000; //  e
         799: data = 8'b00000000; //  f
          //    code x32
         800: data = 8'b00000000; //  0
         801: data = 8'b00000000; //  1
         802: data = 8'b01111100; //  2  *****
         803: data = 8'b11000110; //  3 **   **
         804: data = 8'b00000110; //  4      **
         805: data = 8'b00001100; //  5     **
         806: data = 8'b00011000; //  6    **
         807: data = 8'b00110000; //  7   **
         808: data = 8'b01100000; //  8  **
         809: data = 8'b11000000; //  9 **
         810: data = 8'b11000110; //  a **   **
         811: data = 8'b11111110; //  b *******
         812: data = 8'b00000000; //  c
         813: data = 8'b00000000; //  d
         814: data = 8'b00000000; //  e
         815: data = 8'b00000000; //  f
          //    code x33
         816: data = 8'b00000000; //  0
         817: data = 8'b00000000; //  1
         818: data = 8'b01111100; //  2  *****
         819: data = 8'b11000110; //  3 **   **
         820: data = 8'b00000110; //  4      **
         821: data = 8'b00000110; //  5      **
         822: data = 8'b00111100; //  6   ****
         823: data = 8'b00000110; //  7      **
         824: data = 8'b00000110; //  8      **
         825: data = 8'b00000110; //  9      **
         826: data = 8'b11000110; //  a **   **
         827: data = 8'b01111100; //  b  *****
         828: data = 8'b00000000; //  c
         829: data = 8'b00000000; //  d
         830: data = 8'b00000000; //  e
         831: data = 8'b00000000; //  f
          //    code x34
         832: data = 8'b00000000; //  0
         833: data = 8'b00000000; //  1
         834: data = 8'b00001100; //  2     **
         835: data = 8'b00011100; //  3    ***
         836: data = 8'b00111100; //  4   ****
         837: data = 8'b01101100; //  5  ** **
         838: data = 8'b11001100; //  6 **  **
         839: data = 8'b11111110; //  7 *******
         840: data = 8'b00001100; //  8     **
         841: data = 8'b00001100; //  9     **
         842: data = 8'b00001100; //  a     **
         843: data = 8'b00011110; //  b    ****
         844: data = 8'b00000000; //  c
         845: data = 8'b00000000; //  d
         846: data = 8'b00000000; //  e
         847: data = 8'b00000000; //  f
          //    code x35
         848: data = 8'b00000000; //  0
         849: data = 8'b00000000; //  1
         850: data = 8'b11111110; //  2 *******
         851: data = 8'b11000000; //  3 **
         852: data = 8'b11000000; //  4 **
         853: data = 8'b11000000; //  5 **
         854: data = 8'b11111100; //  6 ******
         855: data = 8'b00000110; //  7      **
         856: data = 8'b00000110; //  8      **
         857: data = 8'b00000110; //  9      **
         858: data = 8'b11000110; //  a **   **
         859: data = 8'b01111100; //  b  *****
         860: data = 8'b00000000; //  c
         861: data = 8'b00000000; //  d
         862: data = 8'b00000000; //  e
         863: data = 8'b00000000; //  f
          //    code x36
         864: data = 8'b00000000; //  0
         865: data = 8'b00000000; //  1
         866: data = 8'b00111000; //  2   ***
         867: data = 8'b01100000; //  3  **
         868: data = 8'b11000000; //  4 **
         869: data = 8'b11000000; //  5 **
         870: data = 8'b11111100; //  6 ******
         871: data = 8'b11000110; //  7 **   **
         872: data = 8'b11000110; //  8 **   **
         873: data = 8'b11000110; //  9 **   **
         874: data = 8'b11000110; //  a **   **
         875: data = 8'b01111100; //  b  *****
         876: data = 8'b00000000; //  c
         877: data = 8'b00000000; //  d
         878: data = 8'b00000000; //  e
         879: data = 8'b00000000; //  f
          //    code x37
         880: data = 8'b00000000; //  0
         881: data = 8'b00000000; //  1
         882: data = 8'b11111110; //  2 *******
         883: data = 8'b11000110; //  3 **   **
         884: data = 8'b00000110; //  4      **
         885: data = 8'b00000110; //  5      **
         886: data = 8'b00001100; //  6     **
         887: data = 8'b00011000; //  7    **
         888: data = 8'b00110000; //  8   **
         889: data = 8'b00110000; //  9   **
         890: data = 8'b00110000; //  a   **
         891: data = 8'b00110000; //  b   **
         892: data = 8'b00000000; //  c
         893: data = 8'b00000000; //  d
         894: data = 8'b00000000; //  e
         895: data = 8'b00000000; //  f
          //    code x38
         896: data = 8'b00000000; //  0
         897: data = 8'b00000000; //  1
         898: data = 8'b01111100; //  2  *****
         899: data = 8'b11000110; //  3 **   **
         900: data = 8'b11000110; //  4 **   **
         901: data = 8'b11000110; //  5 **   **
         902: data = 8'b01111100; //  6  *****
         903: data = 8'b11000110; //  7 **   **
         904: data = 8'b11000110; //  8 **   **
         905: data = 8'b11000110; //  9 **   **
         906: data = 8'b11000110; //  a **   **
         907: data = 8'b01111100; //  b  *****
         908: data = 8'b00000000; //  c
         909: data = 8'b00000000; //  d
         910: data = 8'b00000000; //  e
         911: data = 8'b00000000; //  f
          //    code x39
         912: data = 8'b00000000; //  0
         913: data = 8'b00000000; //  1
         914: data = 8'b01111100; //  2  *****
         915: data = 8'b11000110; //  3 **   **
         916: data = 8'b11000110; //  4 **   **
         917: data = 8'b11000110; //  5 **   **
         918: data = 8'b01111110; //  6  ******
         919: data = 8'b00000110; //  7      **
         920: data = 8'b00000110; //  8      **
         921: data = 8'b00000110; //  9      **
         922: data = 8'b00001100; //  a     **
         923: data = 8'b01111000; //  b  ****
         924: data = 8'b00000000; //  c
         925: data = 8'b00000000; //  d
         926: data = 8'b00000000; //  e
         927: data = 8'b00000000; //  f
          //    code x3a
         928: data = 8'b00000000; //  0
         929: data = 8'b00000000; //  1
         930: data = 8'b00000000; //  2
         931: data = 8'b00000000; //  3
         932: data = 8'b00011000; //  4    **
         933: data = 8'b00011000; //  5    **
         934: data = 8'b00000000; //  6
         935: data = 8'b00000000; //  7
         936: data = 8'b00000000; //  8
         937: data = 8'b00011000; //  9    **
         938: data = 8'b00011000; //  a    **
         939: data = 8'b00000000; //  b
         940: data = 8'b00000000; //  c
         941: data = 8'b00000000; //  d
         942: data = 8'b00000000; //  e
         943: data = 8'b00000000; //  f
          //    code x3b
         944: data = 8'b00000000; //  0
         945: data = 8'b00000000; //  1
         946: data = 8'b00000000; //  2
         947: data = 8'b00000000; //  3
         948: data = 8'b00011000; //  4    **
         949: data = 8'b00011000; //  5    **
         950: data = 8'b00000000; //  6
         951: data = 8'b00000000; //  7
         952: data = 8'b00000000; //  8
         953: data = 8'b00011000; //  9    **
         954: data = 8'b00011000; //  a    **
         955: data = 8'b00110000; //  b   **
         956: data = 8'b00000000; //  c
         957: data = 8'b00000000; //  d
         958: data = 8'b00000000; //  e
         959: data = 8'b00000000; //  f
          //    code x3c
         960: data = 8'b00000000; //  0
         961: data = 8'b00000000; //  1
         962: data = 8'b00000000; //  2
         963: data = 8'b00000110; //  3      **
         964: data = 8'b00001100; //  4     **
         965: data = 8'b00011000; //  5    **
         966: data = 8'b00110000; //  6   **
         967: data = 8'b01100000; //  7  **
         968: data = 8'b00110000; //  8   **
         969: data = 8'b00011000; //  9    **
         970: data = 8'b00001100; //  a     **
         971: data = 8'b00000110; //  b      **
         972: data = 8'b00000000; //  c
         973: data = 8'b00000000; //  d
         974: data = 8'b00000000; //  e
         975: data = 8'b00000000; //  f
          //    code x3d
         976: data = 8'b00000000; //  0
         977: data = 8'b00000000; //  1
         978: data = 8'b00000000; //  2
         979: data = 8'b00000000; //  3
         980: data = 8'b00000000; //  4
         981: data = 8'b01111110; //  5  ******
         982: data = 8'b00000000; //  6
         983: data = 8'b00000000; //  7
         984: data = 8'b01111110; //  8  ******
         985: data = 8'b00000000; //  9
         986: data = 8'b00000000; //  a
         987: data = 8'b00000000; //  b
         988: data = 8'b00000000; //  c
         989: data = 8'b00000000; //  d
         990: data = 8'b00000000; //  e
         991: data = 8'b00000000; //  f
          //    code x3e
         992: data = 8'b00000000; //  0
         993: data = 8'b00000000; //  1
         994: data = 8'b00000000; //  2
         995: data = 8'b01100000; //  3  **
         996: data = 8'b00110000; //  4   **
         997: data = 8'b00011000; //  5    **
         998: data = 8'b00001100; //  6     **
         999: data = 8'b00000110; //  7      **
        1000: data = 8'b00001100; //  8     **
        1001: data = 8'b00011000; //  9    **
        1002: data = 8'b00110000; //  a   **
        1003: data = 8'b01100000; //  b  **
        1004: data = 8'b00000000; //  c
        1005: data = 8'b00000000; //  d
        1006: data = 8'b00000000; //  e
        1007: data = 8'b00000000; //  f
          //    code x3f
        1008: data = 8'b00000000; //  0
        1009: data = 8'b00000000; //  1
        1010: data = 8'b01111100; //  2  *****
        1011: data = 8'b11000110; //  3 **   **
        1012: data = 8'b11000110; //  4 **   **
        1013: data = 8'b00001100; //  5     **
        1014: data = 8'b00011000; //  6    **
        1015: data = 8'b00011000; //  7    **
        1016: data = 8'b00011000; //  8    **
        1017: data = 8'b00000000; //  9
        1018: data = 8'b00011000; //  a    **
        1019: data = 8'b00011000; //  b    **
        1020: data = 8'b00000000; //  c
        1021: data = 8'b00000000; //  d
        1022: data = 8'b00000000; //  e
        1023: data = 8'b00000000; //  f
          //    code x40
        1024: data = 8'b00000000; //  0
        1025: data = 8'b00000000; //  1
        1026: data = 8'b01111100; //  2  *****
        1027: data = 8'b11000110; //  3 **   **
        1028: data = 8'b11000110; //  4 **   **
        1029: data = 8'b11000110; //  5 **   **
        1030: data = 8'b11011110; //  6 ** ****
        1031: data = 8'b11011110; //  7 ** ****
        1032: data = 8'b11011110; //  8 ** ****
        1033: data = 8'b11011100; //  9 ** ***
        1034: data = 8'b11000000; //  a **
        1035: data = 8'b01111100; //  b  *****
        1036: data = 8'b00000000; //  c
        1037: data = 8'b00000000; //  d
        1038: data = 8'b00000000; //  e
        1039: data = 8'b00000000; //  f
          //    code x41
        1040: data = 8'b00000000; //  0
        1041: data = 8'b00000000; //  1
        1042: data = 8'b00010000; //  2    *
        1043: data = 8'b00111000; //  3   ***
        1044: data = 8'b01101100; //  4  ** **
        1045: data = 8'b11000110; //  5 **   **
        1046: data = 8'b11000110; //  6 **   **
        1047: data = 8'b11111110; //  7 *******
        1048: data = 8'b11000110; //  8 **   **
        1049: data = 8'b11000110; //  9 **   **
        1050: data = 8'b11000110; //  a **   **
        1051: data = 8'b11000110; //  b **   **
        1052: data = 8'b00000000; //  c
        1053: data = 8'b00000000; //  d
        1054: data = 8'b00000000; //  e
        1055: data = 8'b00000000; //  f
          //    code x42
        1056: data = 8'b00000000; //  0
        1057: data = 8'b00000000; //  1
        1058: data = 8'b11111100; //  2 ******
        1059: data = 8'b01100110; //  3  **  **
        1060: data = 8'b01100110; //  4  **  **
        1061: data = 8'b01100110; //  5  **  **
        1062: data = 8'b01111100; //  6  *****
        1063: data = 8'b01100110; //  7  **  **
        1064: data = 8'b01100110; //  8  **  **
        1065: data = 8'b01100110; //  9  **  **
        1066: data = 8'b01100110; //  a  **  **
        1067: data = 8'b11111100; //  b ******
        1068: data = 8'b00000000; //  c
        1069: data = 8'b00000000; //  d
        1070: data = 8'b00000000; //  e
        1071: data = 8'b00000000; //  f
          //    code x43
        1072: data = 8'b00000000; //  0
        1073: data = 8'b00000000; //  1
        1074: data = 8'b00111100; //  2   ****
        1075: data = 8'b01100110; //  3  **  **
        1076: data = 8'b11000010; //  4 **    *
        1077: data = 8'b11000000; //  5 **
        1078: data = 8'b11000000; //  6 **
        1079: data = 8'b11000000; //  7 **
        1080: data = 8'b11000000; //  8 **
        1081: data = 8'b11000010; //  9 **    *
        1082: data = 8'b01100110; //  a  **  **
        1083: data = 8'b00111100; //  b   ****
        1084: data = 8'b00000000; //  c
        1085: data = 8'b00000000; //  d
        1086: data = 8'b00000000; //  e
        1087: data = 8'b00000000; //  f
          //    code x44
        1088: data = 8'b00000000; //  0
        1089: data = 8'b00000000; //  1
        1090: data = 8'b11111000; //  2 *****
        1091: data = 8'b01101100; //  3  ** **
        1092: data = 8'b01100110; //  4  **  **
        1093: data = 8'b01100110; //  5  **  **
        1094: data = 8'b01100110; //  6  **  **
        1095: data = 8'b01100110; //  7  **  **
        1096: data = 8'b01100110; //  8  **  **
        1097: data = 8'b01100110; //  9  **  **
        1098: data = 8'b01101100; //  a  ** **
        1099: data = 8'b11111000; //  b *****
        1100: data = 8'b00000000; //  c
        1101: data = 8'b00000000; //  d
        1102: data = 8'b00000000; //  e
        1103: data = 8'b00000000; //  f
          //    code x45
        1104: data = 8'b00000000; //  0
        1105: data = 8'b00000000; //  1
        1106: data = 8'b11111110; //  2 *******
        1107: data = 8'b01100110; //  3  **  **
        1108: data = 8'b01100010; //  4  **   *
        1109: data = 8'b01101000; //  5  ** *
        1110: data = 8'b01111000; //  6  ****
        1111: data = 8'b01101000; //  7  ** *
        1112: data = 8'b01100000; //  8  **
        1113: data = 8'b01100010; //  9  **   *
        1114: data = 8'b01100110; //  a  **  **
        1115: data = 8'b11111110; //  b *******
        1116: data = 8'b00000000; //  c
        1117: data = 8'b00000000; //  d
        1118: data = 8'b00000000; //  e
        1119: data = 8'b00000000; //  f
          //    code x46
        1120: data = 8'b00000000; //  0
        1121: data = 8'b00000000; //  1
        1122: data = 8'b11111110; //  2 *******
        1123: data = 8'b01100110; //  3  **  **
        1124: data = 8'b01100010; //  4  **   *
        1125: data = 8'b01101000; //  5  ** *
        1126: data = 8'b01111000; //  6  ****
        1127: data = 8'b01101000; //  7  ** *
        1128: data = 8'b01100000; //  8  **
        1129: data = 8'b01100000; //  9  **
        1130: data = 8'b01100000; //  a  **
        1131: data = 8'b11110000; //  b ****
        1132: data = 8'b00000000; //  c
        1133: data = 8'b00000000; //  d
        1134: data = 8'b00000000; //  e
        1135: data = 8'b00000000; //  f
          //    code x47
        1136: data = 8'b00000000; //  0
        1137: data = 8'b00000000; //  1
        1138: data = 8'b00111100; //  2   ****
        1139: data = 8'b01100110; //  3  **  **
        1140: data = 8'b11000010; //  4 **    *
        1141: data = 8'b11000000; //  5 **
        1142: data = 8'b11000000; //  6 **
        1143: data = 8'b11011110; //  7 ** ****
        1144: data = 8'b11000110; //  8 **   **
        1145: data = 8'b11000110; //  9 **   **
        1146: data = 8'b01100110; //  a  **  **
        1147: data = 8'b00111010; //  b   *** *
        1148: data = 8'b00000000; //  c
        1149: data = 8'b00000000; //  d
        1150: data = 8'b00000000; //  e
        1151: data = 8'b00000000; //  f
          //    code x48
        1152: data = 8'b00000000; //  0
        1153: data = 8'b00000000; //  1
        1154: data = 8'b11000110; //  2 **   **
        1155: data = 8'b11000110; //  3 **   **
        1156: data = 8'b11000110; //  4 **   **
        1157: data = 8'b11000110; //  5 **   **
        1158: data = 8'b11111110; //  6 *******
        1159: data = 8'b11000110; //  7 **   **
        1160: data = 8'b11000110; //  8 **   **
        1161: data = 8'b11000110; //  9 **   **
        1162: data = 8'b11000110; //  a **   **
        1163: data = 8'b11000110; //  b **   **
        1164: data = 8'b00000000; //  c
        1165: data = 8'b00000000; //  d
        1166: data = 8'b00000000; //  e
        1167: data = 8'b00000000; //  f
          //    code x49
        1168: data = 8'b00000000; //  0
        1169: data = 8'b00000000; //  1
        1170: data = 8'b00111100; //  2   ****
        1171: data = 8'b00011000; //  3    **
        1172: data = 8'b00011000; //  4    **
        1173: data = 8'b00011000; //  5    **
        1174: data = 8'b00011000; //  6    **
        1175: data = 8'b00011000; //  7    **
        1176: data = 8'b00011000; //  8    **
        1177: data = 8'b00011000; //  9    **
        1178: data = 8'b00011000; //  a    **
        1179: data = 8'b00111100; //  b   ****
        1180: data = 8'b00000000; //  c
        1181: data = 8'b00000000; //  d
        1182: data = 8'b00000000; //  e
        1183: data = 8'b00000000; //  f
          //    code x4a
        1184: data = 8'b00000000; //  0
        1185: data = 8'b00000000; //  1
        1186: data = 8'b00011110; //  2    ****
        1187: data = 8'b00001100; //  3     **
        1188: data = 8'b00001100; //  4     **
        1189: data = 8'b00001100; //  5     **
        1190: data = 8'b00001100; //  6     **
        1191: data = 8'b00001100; //  7     **
        1192: data = 8'b11001100; //  8 **  **
        1193: data = 8'b11001100; //  9 **  **
        1194: data = 8'b11001100; //  a **  **
        1195: data = 8'b01111000; //  b  ****
        1196: data = 8'b00000000; //  c
        1197: data = 8'b00000000; //  d
        1198: data = 8'b00000000; //  e
        1199: data = 8'b00000000; //  f
          //    code x4b
        1200: data = 8'b00000000; //  0
        1201: data = 8'b00000000; //  1
        1202: data = 8'b11100110; //  2 ***  **
        1203: data = 8'b01100110; //  3  **  **
        1204: data = 8'b01100110; //  4  **  **
        1205: data = 8'b01101100; //  5  ** **
        1206: data = 8'b01111000; //  6  ****
        1207: data = 8'b01111000; //  7  ****
        1208: data = 8'b01101100; //  8  ** **
        1209: data = 8'b01100110; //  9  **  **
        1210: data = 8'b01100110; //  a  **  **
        1211: data = 8'b11100110; //  b ***  **
        1212: data = 8'b00000000; //  c
        1213: data = 8'b00000000; //  d
        1214: data = 8'b00000000; //  e
        1215: data = 8'b00000000; //  f
          //    code x4c
        1216: data = 8'b00000000; //  0
        1217: data = 8'b00000000; //  1
        1218: data = 8'b11110000; //  2 ****
        1219: data = 8'b01100000; //  3  **
        1220: data = 8'b01100000; //  4  **
        1221: data = 8'b01100000; //  5  **
        1222: data = 8'b01100000; //  6  **
        1223: data = 8'b01100000; //  7  **
        1224: data = 8'b01100000; //  8  **
        1225: data = 8'b01100010; //  9  **   *
        1226: data = 8'b01100110; //  a  **  **
        1227: data = 8'b11111110; //  b *******
        1228: data = 8'b00000000; //  c
        1229: data = 8'b00000000; //  d
        1230: data = 8'b00000000; //  e
        1231: data = 8'b00000000; //  f
          //    code x4d
        1232: data = 8'b00000000; //  0
        1233: data = 8'b00000000; //  1
        1234: data = 8'b11000011; //  2 **    **
        1235: data = 8'b11100111; //  3 ***  ***
        1236: data = 8'b11111111; //  4 ********
        1237: data = 8'b11111111; //  5 ********
        1238: data = 8'b11011011; //  6 ** ** **
        1239: data = 8'b11000011; //  7 **    **
        1240: data = 8'b11000011; //  8 **    **
        1241: data = 8'b11000011; //  9 **    **
        1242: data = 8'b11000011; //  a **    **
        1243: data = 8'b11000011; //  b **    **
        1244: data = 8'b00000000; //  c
        1245: data = 8'b00000000; //  d
        1246: data = 8'b00000000; //  e
        1247: data = 8'b00000000; //  f
          //    code x4e
        1248: data = 8'b00000000; //  0
        1249: data = 8'b00000000; //  1
        1250: data = 8'b11000110; //  2 **   **
        1251: data = 8'b11100110; //  3 ***  **
        1252: data = 8'b11110110; //  4 **** **
        1253: data = 8'b11111110; //  5 *******
        1254: data = 8'b11011110; //  6 ** ****
        1255: data = 8'b11001110; //  7 **  ***
        1256: data = 8'b11000110; //  8 **   **
        1257: data = 8'b11000110; //  9 **   **
        1258: data = 8'b11000110; //  a **   **
        1259: data = 8'b11000110; //  b **   **
        1260: data = 8'b00000000; //  c
        1261: data = 8'b00000000; //  d
        1262: data = 8'b00000000; //  e
        1263: data = 8'b00000000; //  f
          //    code x4f
        1264: data = 8'b00000000; //  0
        1265: data = 8'b00000000; //  1
        1266: data = 8'b01111100; //  2  *****
        1267: data = 8'b11000110; //  3 **   **
        1268: data = 8'b11000110; //  4 **   **
        1269: data = 8'b11000110; //  5 **   **
        1270: data = 8'b11000110; //  6 **   **
        1271: data = 8'b11000110; //  7 **   **
        1272: data = 8'b11000110; //  8 **   **
        1273: data = 8'b11000110; //  9 **   **
        1274: data = 8'b11000110; //  a **   **
        1275: data = 8'b01111100; //  b  *****
        1276: data = 8'b00000000; //  c
        1277: data = 8'b00000000; //  d
        1278: data = 8'b00000000; //  e
        1279: data = 8'b00000000; //  f
          //    code x50
        1280: data = 8'b00000000; //  0
        1281: data = 8'b00000000; //  1
        1282: data = 8'b11111100; //  2 ******
        1283: data = 8'b01100110; //  3  **  **
        1284: data = 8'b01100110; //  4  **  **
        1285: data = 8'b01100110; //  5  **  **
        1286: data = 8'b01111100; //  6  *****
        1287: data = 8'b01100000; //  7  **
        1288: data = 8'b01100000; //  8  **
        1289: data = 8'b01100000; //  9  **
        1290: data = 8'b01100000; //  a  **
        1291: data = 8'b11110000; //  b ****
        1292: data = 8'b00000000; //  c
        1293: data = 8'b00000000; //  d
        1294: data = 8'b00000000; //  e
        1295: data = 8'b00000000; //  f
          //    code x510
        1296: data = 8'b00000000; //  0
        1297: data = 8'b00000000; //  1
        1298: data = 8'b01111100; //  2  *****
        1299: data = 8'b11000110; //  3 **   **
        1300: data = 8'b11000110; //  4 **   **
        1301: data = 8'b11000110; //  5 **   **
        1302: data = 8'b11000110; //  6 **   **
        1303: data = 8'b11000110; //  7 **   **
        1304: data = 8'b11000110; //  8 **   **
        1305: data = 8'b11010110; //  9 ** * **
        1306: data = 8'b11011110; //  a ** ****
        1307: data = 8'b01111100; //  b  *****
        1308: data = 8'b00001100; //  c     **
        1309: data = 8'b00001110; //  d     ***
        1310: data = 8'b00000000; //  e
        1311: data = 8'b00000000; //  f
          //    code x52
        1312: data = 8'b00000000; //  0
        1313: data = 8'b00000000; //  1
        1314: data = 8'b11111100; //  2 ******
        1315: data = 8'b01100110; //  3  **  **
        1316: data = 8'b01100110; //  4  **  **
        1317: data = 8'b01100110; //  5  **  **
        1318: data = 8'b01111100; //  6  *****
        1319: data = 8'b01101100; //  7  ** **
        1320: data = 8'b01100110; //  8  **  **
        1321: data = 8'b01100110; //  9  **  **
        1322: data = 8'b01100110; //  a  **  **
        1323: data = 8'b11100110; //  b ***  **
        1324: data = 8'b00000000; //  c
        1325: data = 8'b00000000; //  d
        1326: data = 8'b00000000; //  e
        1327: data = 8'b00000000; //  f
          //    code x53
        1328: data = 8'b00000000; //  0
        1329: data = 8'b00000000; //  1
        1330: data = 8'b01111100; //  2  *****
        1331: data = 8'b11000110; //  3 **   **
        1332: data = 8'b11000110; //  4 **   **
        1333: data = 8'b01100000; //  5  **
        1334: data = 8'b00111000; //  6   ***
        1335: data = 8'b00001100; //  7     **
        1336: data = 8'b00000110; //  8      **
        1337: data = 8'b11000110; //  9 **   **
        1338: data = 8'b11000110; //  a **   **
        1339: data = 8'b01111100; //  b  *****
        1340: data = 8'b00000000; //  c
        1341: data = 8'b00000000; //  d
        1342: data = 8'b00000000; //  e
        1343: data = 8'b00000000; //  f
          //    code x54
        1344: data = 8'b00000000; //  0
        1345: data = 8'b00000000; //  1
        1346: data = 8'b11111111; //  2 ********
        1347: data = 8'b11011011; //  3 ** ** **
        1348: data = 8'b10011001; //  4 *  **  *
        1349: data = 8'b00011000; //  5    **
        1350: data = 8'b00011000; //  6    **
        1351: data = 8'b00011000; //  7    **
        1352: data = 8'b00011000; //  8    **
        1353: data = 8'b00011000; //  9    **
        1354: data = 8'b00011000; //  a    **
        1355: data = 8'b00111100; //  b   ****
        1356: data = 8'b00000000; //  c
        1357: data = 8'b00000000; //  d
        1358: data = 8'b00000000; //  e
        1359: data = 8'b00000000; //  f
          //    code x55
        1360: data = 8'b00000000; //  0
        1361: data = 8'b00000000; //  1
        1362: data = 8'b11000110; //  2 **   **
        1363: data = 8'b11000110; //  3 **   **
        1364: data = 8'b11000110; //  4 **   **
        1365: data = 8'b11000110; //  5 **   **
        1366: data = 8'b11000110; //  6 **   **
        1367: data = 8'b11000110; //  7 **   **
        1368: data = 8'b11000110; //  8 **   **
        1369: data = 8'b11000110; //  9 **   **
        1370: data = 8'b11000110; //  a **   **
        1371: data = 8'b01111100; //  b  *****
        1372: data = 8'b00000000; //  c
        1373: data = 8'b00000000; //  d
        1374: data = 8'b00000000; //  e
        1375: data = 8'b00000000; //  f
          //    code x56
        1376: data = 8'b00000000; //  0
        1377: data = 8'b00000000; //  1
        1378: data = 8'b11000011; //  2 **    **
        1379: data = 8'b11000011; //  3 **    **
        1380: data = 8'b11000011; //  4 **    **
        1381: data = 8'b11000011; //  5 **    **
        1382: data = 8'b11000011; //  6 **    **
        1383: data = 8'b11000011; //  7 **    **
        1384: data = 8'b11000011; //  8 **    **
        1385: data = 8'b01100110; //  9  **  **
        1386: data = 8'b00111100; //  a   ****
        1387: data = 8'b00011000; //  b    **
        1388: data = 8'b00000000; //  c
        1389: data = 8'b00000000; //  d
        1390: data = 8'b00000000; //  e
        1391: data = 8'b00000000; //  f
          //    code x57
        1392: data = 8'b00000000; //  0
        1393: data = 8'b00000000; //  1
        1394: data = 8'b11000011; //  2 **    **
        1395: data = 8'b11000011; //  3 **    **
        1396: data = 8'b11000011; //  4 **    **
        1397: data = 8'b11000011; //  5 **    **
        1398: data = 8'b11000011; //  6 **    **
        1399: data = 8'b11011011; //  7 ** ** **
        1400: data = 8'b11011011; //  8 ** ** **
        1401: data = 8'b11111111; //  9 ********
        1402: data = 8'b01100110; //  a  **  **
        1403: data = 8'b01100110; //  b  **  **
        1404: data = 8'b00000000; //  c
        1405: data = 8'b00000000; //  d
        1406: data = 8'b00000000; //  e
        1407: data = 8'b00000000; //  f
          //    code x58
        1408: data = 8'b00000000; //  0
        1409: data = 8'b00000000; //  1
        1410: data = 8'b11000011; //  2 **    **
        1411: data = 8'b11000011; //  3 **    **
        1412: data = 8'b01100110; //  4  **  **
        1413: data = 8'b00111100; //  5   ****
        1414: data = 8'b00011000; //  6    **
        1415: data = 8'b00011000; //  7    **
        1416: data = 8'b00111100; //  8   ****
        1417: data = 8'b01100110; //  9  **  **
        1418: data = 8'b11000011; //  a **    **
        1419: data = 8'b11000011; //  b **    **
        1420: data = 8'b00000000; //  c
        1421: data = 8'b00000000; //  d
        1422: data = 8'b00000000; //  e
        1423: data = 8'b00000000; //  f
          //    code x59
        1424: data = 8'b00000000; //  0
        1425: data = 8'b00000000; //  1
        1426: data = 8'b11000011; //  2 **    **
        1427: data = 8'b11000011; //  3 **    **
        1428: data = 8'b11000011; //  4 **    **
        1429: data = 8'b01100110; //  5  **  **
        1430: data = 8'b00111100; //  6   ****
        1431: data = 8'b00011000; //  7    **
        1432: data = 8'b00011000; //  8    **
        1433: data = 8'b00011000; //  9    **
        1434: data = 8'b00011000; //  a    **
        1435: data = 8'b00111100; //  b   ****
        1436: data = 8'b00000000; //  c
        1437: data = 8'b00000000; //  d
        1438: data = 8'b00000000; //  e
        1439: data = 8'b00000000; //  f
          //    code x5a
        1440: data = 8'b00000000; //  0
        1441: data = 8'b00000000; //  1
        1442: data = 8'b11111111; //  2 ********
        1443: data = 8'b11000011; //  3 **    **
        1444: data = 8'b10000110; //  4 *    **
        1445: data = 8'b00001100; //  5     **
        1446: data = 8'b00011000; //  6    **
        1447: data = 8'b00110000; //  7   **
        1448: data = 8'b01100000; //  8  **
        1449: data = 8'b11000001; //  9 **     *
        1450: data = 8'b11000011; //  a **    **
        1451: data = 8'b11111111; //  b ********
        1452: data = 8'b00000000; //  c
        1453: data = 8'b00000000; //  d
        1454: data = 8'b00000000; //  e
        1455: data = 8'b00000000; //  f
          //    code x5b
        1456: data = 8'b00000000; //  0
        1457: data = 8'b00000000; //  1
        1458: data = 8'b00111100; //  2   ****
        1459: data = 8'b00110000; //  3   **
        1460: data = 8'b00110000; //  4   **
        1461: data = 8'b00110000; //  5   **
        1462: data = 8'b00110000; //  6   **
        1463: data = 8'b00110000; //  7   **
        1464: data = 8'b00110000; //  8   **
        1465: data = 8'b00110000; //  9   **
        1466: data = 8'b00110000; //  a   **
        1467: data = 8'b00111100; //  b   ****
        1468: data = 8'b00000000; //  c
        1469: data = 8'b00000000; //  d
        1470: data = 8'b00000000; //  e
        1471: data = 8'b00000000; //  f
          //    code x5c
        1472: data = 8'b00000000; //  0
        1473: data = 8'b00000000; //  1
        1474: data = 8'b00000000; //  2
        1475: data = 8'b10000000; //  3 *
        1476: data = 8'b11000000; //  4 **
        1477: data = 8'b11100000; //  5 ***
        1478: data = 8'b01110000; //  6  ***
        1479: data = 8'b00111000; //  7   ***
        1480: data = 8'b00011100; //  8    ***
        1481: data = 8'b00001110; //  9     ***
        1482: data = 8'b00000110; //  a      **
        1483: data = 8'b00000010; //  b       *
        1484: data = 8'b00000000; //  c
        1485: data = 8'b00000000; //  d
        1486: data = 8'b00000000; //  e
        1487: data = 8'b00000000; //  f
          //    code x5d
        1488: data = 8'b00000000; //  0
        1489: data = 8'b00000000; //  1
        1490: data = 8'b00111100; //  2   ****
        1491: data = 8'b00001100; //  3     **
        1492: data = 8'b00001100; //  4     **
        1493: data = 8'b00001100; //  5     **
        1494: data = 8'b00001100; //  6     **
        1495: data = 8'b00001100; //  7     **
        1496: data = 8'b00001100; //  8     **
        1497: data = 8'b00001100; //  9     **
        1498: data = 8'b00001100; //  a     **
        1499: data = 8'b00111100; //  b   ****
        1500: data = 8'b00000000; //  c
        1501: data = 8'b00000000; //  d
        1502: data = 8'b00000000; //  e
        1503: data = 8'b00000000; //  f
          //    code x5e
        1504: data = 8'b00010000; //  0    *
        1505: data = 8'b00111000; //  1   ***
        1506: data = 8'b01101100; //  2  ** **
        1507: data = 8'b11000110; //  3 **   **
        1508: data = 8'b00000000; //  4
        1509: data = 8'b00000000; //  5
        1510: data = 8'b00000000; //  6
        1511: data = 8'b00000000; //  7
        1512: data = 8'b00000000; //  8
        1513: data = 8'b00000000; //  9
        1514: data = 8'b00000000; //  a
        1515: data = 8'b00000000; //  b
        1516: data = 8'b00000000; //  c
        1517: data = 8'b00000000; //  d
        1518: data = 8'b00000000; //  e
        1519: data = 8'b00000000; //  f
          //    code x5f
        1520: data = 8'b00000000; //  0
        1521: data = 8'b00000000; //  1
        1522: data = 8'b00000000; //  2
        1523: data = 8'b00000000; //  3
        1524: data = 8'b00000000; //  4
        1525: data = 8'b00000000; //  5
        1526: data = 8'b00000000; //  6
        1527: data = 8'b00000000; //  7
        1528: data = 8'b00000000; //  8
        1529: data = 8'b00000000; //  9
        1530: data = 8'b00000000; //  a
        1531: data = 8'b00000000; //  b
        1532: data = 8'b00000000; //  c
        1533: data = 8'b11111111; //  d ********
        1534: data = 8'b00000000; //  e
        1535: data = 8'b00000000; //  f
          //    code x60
        1536: data = 8'b00110000; //  0   **
        1537: data = 8'b00110000; //  1   **
        1538: data = 8'b00011000; //  2    **
        1539: data = 8'b00000000; //  3
        1540: data = 8'b00000000; //  4
        1541: data = 8'b00000000; //  5
        1542: data = 8'b00000000; //  6
        1543: data = 8'b00000000; //  7
        1544: data = 8'b00000000; //  8
        1545: data = 8'b00000000; //  9
        1546: data = 8'b00000000; //  a
        1547: data = 8'b00000000; //  b
        1548: data = 8'b00000000; //  c
        1549: data = 8'b00000000; //  d
        1550: data = 8'b00000000; //  e
        1551: data = 8'b00000000; //  f
          //    code x61
        1552: data = 8'b00000000; //  0
        1553: data = 8'b00000000; //  1
        1554: data = 8'b00000000; //  2
        1555: data = 8'b00000000; //  3
        1556: data = 8'b00000000; //  4
        1557: data = 8'b01111000; //  5  ****
        1558: data = 8'b00001100; //  6     **
        1559: data = 8'b01111100; //  7  *****
        1560: data = 8'b11001100; //  8 **  **
        1561: data = 8'b11001100; //  9 **  **
        1562: data = 8'b11001100; //  a **  **
        1563: data = 8'b01110110; //  b  *** **
        1564: data = 8'b00000000; //  c
        1565: data = 8'b00000000; //  d
        1566: data = 8'b00000000; //  e
        1567: data = 8'b00000000; //  f
          //    code x62
        1568: data = 8'b00000000; //  0
        1569: data = 8'b00000000; //  1
        1570: data = 8'b11100000; //  2  ***
        1571: data = 8'b01100000; //  3   **
        1572: data = 8'b01100000; //  4   **
        1573: data = 8'b01111000; //  5   ****
        1574: data = 8'b01101100; //  6   ** **
        1575: data = 8'b01100110; //  7   **  **
        1576: data = 8'b01100110; //  8   **  **
        1577: data = 8'b01100110; //  9   **  **
        1578: data = 8'b01100110; //  a   **  **
        1579: data = 8'b01111100; //  b   *****
        1580: data = 8'b00000000; //  c
        1581: data = 8'b00000000; //  d
        1582: data = 8'b00000000; //  e
        1583: data = 8'b00000000; //  f
          //    code x63
        1584: data = 8'b00000000; //  0
        1585: data = 8'b00000000; //  1
        1586: data = 8'b00000000; //  2
        1587: data = 8'b00000000; //  3
        1588: data = 8'b00000000; //  4
        1589: data = 8'b01111100; //  5  *****
        1590: data = 8'b11000110; //  6 **   **
        1591: data = 8'b11000000; //  7 **
        1592: data = 8'b11000000; //  8 **
        1593: data = 8'b11000000; //  9 **
        1594: data = 8'b11000110; //  a **   **
        1595: data = 8'b01111100; //  b  *****
        1596: data = 8'b00000000; //  c
        1597: data = 8'b00000000; //  d
        1598: data = 8'b00000000; //  e
        1599: data = 8'b00000000; //  f
          //    code x64
        1600: data = 8'b00000000; //  0
        1601: data = 8'b00000000; //  1
        1602: data = 8'b00011100; //  2    ***
        1603: data = 8'b00001100; //  3     **
        1604: data = 8'b00001100; //  4     **
        1605: data = 8'b00111100; //  5   ****
        1606: data = 8'b01101100; //  6  ** **
        1607: data = 8'b11001100; //  7 **  **
        1608: data = 8'b11001100; //  8 **  **
        1609: data = 8'b11001100; //  9 **  **
        1610: data = 8'b11001100; //  a **  **
        1611: data = 8'b01110110; //  b  *** **
        1612: data = 8'b00000000; //  c
        1613: data = 8'b00000000; //  d
        1614: data = 8'b00000000; //  e
        1615: data = 8'b00000000; //  f
          //    code x65
        1616: data = 8'b00000000; //  0
        1617: data = 8'b00000000; //  1
        1618: data = 8'b00000000; //  2
        1619: data = 8'b00000000; //  3
        1620: data = 8'b00000000; //  4
        1621: data = 8'b01111100; //  5  *****
        1622: data = 8'b11000110; //  6 **   **
        1623: data = 8'b11111110; //  7 *******
        1624: data = 8'b11000000; //  8 **
        1625: data = 8'b11000000; //  9 **
        1626: data = 8'b11000110; //  a **   **
        1627: data = 8'b01111100; //  b  *****
        1628: data = 8'b00000000; //  c
        1629: data = 8'b00000000; //  d
        1630: data = 8'b00000000; //  e
        1631: data = 8'b00000000; //  f
          //    code x66
        1632: data = 8'b00000000; //  0
        1633: data = 8'b00000000; //  1
        1634: data = 8'b00111000; //  2   ***
        1635: data = 8'b01101100; //  3  ** **
        1636: data = 8'b01100100; //  4  **  *
        1637: data = 8'b01100000; //  5  **
        1638: data = 8'b11110000; //  6 ****
        1639: data = 8'b01100000; //  7  **
        1640: data = 8'b01100000; //  8  **
        1641: data = 8'b01100000; //  9  **
        1642: data = 8'b01100000; //  a  **
        1643: data = 8'b11110000; //  b ****
        1644: data = 8'b00000000; //  c
        1645: data = 8'b00000000; //  d
        1646: data = 8'b00000000; //  e
        1647: data = 8'b00000000; //  f
          //    code x67
        1648: data = 8'b00000000; //  0
        1649: data = 8'b00000000; //  1
        1650: data = 8'b00000000; //  2
        1651: data = 8'b00000000; //  3
        1652: data = 8'b00000000; //  4
        1653: data = 8'b01110110; //  5  *** **
        1654: data = 8'b11001100; //  6 **  **
        1655: data = 8'b11001100; //  7 **  **
        1656: data = 8'b11001100; //  8 **  **
        1657: data = 8'b11001100; //  9 **  **
        1658: data = 8'b11001100; //  a **  **
        1659: data = 8'b01111100; //  b  *****
        1660: data = 8'b00001100; //  c     **
        1661: data = 8'b11001100; //  d **  **
        1662: data = 8'b01111000; //  e  ****
        1663: data = 8'b00000000; //  f
          //    code x68
        1664: data = 8'b00000000; //  0
        1665: data = 8'b00000000; //  1
        1666: data = 8'b11100000; //  2 ***
        1667: data = 8'b01100000; //  3  **
        1668: data = 8'b01100000; //  4  **
        1669: data = 8'b01101100; //  5  ** **
        1670: data = 8'b01110110; //  6  *** **
        1671: data = 8'b01100110; //  7  **  **
        1672: data = 8'b01100110; //  8  **  **
        1673: data = 8'b01100110; //  9  **  **
        1674: data = 8'b01100110; //  a  **  **
        1675: data = 8'b11100110; //  b ***  **
        1676: data = 8'b00000000; //  c
        1677: data = 8'b00000000; //  d
        1678: data = 8'b00000000; //  e
        1679: data = 8'b00000000; //  f
          //    code x69
        1680: data = 8'b00000000; //  0
        1681: data = 8'b00000000; //  1
        1682: data = 8'b00011000; //  2    **
        1683: data = 8'b00011000; //  3    **
        1684: data = 8'b00000000; //  4
        1685: data = 8'b00111000; //  5   ***
        1686: data = 8'b00011000; //  6    **
        1687: data = 8'b00011000; //  7    **
        1688: data = 8'b00011000; //  8    **
        1689: data = 8'b00011000; //  9    **
        1690: data = 8'b00011000; //  a    **
        1691: data = 8'b00111100; //  b   ****
        1692: data = 8'b00000000; //  c
        1693: data = 8'b00000000; //  d
        1694: data = 8'b00000000; //  e
        1695: data = 8'b00000000; //  f
          //    code x6a
        1696: data = 8'b00000000; //  0
        1697: data = 8'b00000000; //  1
        1698: data = 8'b00000110; //  2      **
        1699: data = 8'b00000110; //  3      **
        1700: data = 8'b00000000; //  4
        1701: data = 8'b00001110; //  5     ***
        1702: data = 8'b00000110; //  6      **
        1703: data = 8'b00000110; //  7      **
        1704: data = 8'b00000110; //  8      **
        1705: data = 8'b00000110; //  9      **
        1706: data = 8'b00000110; //  a      **
        1707: data = 8'b00000110; //  b      **
        1708: data = 8'b01100110; //  c  **  **
        1709: data = 8'b01100110; //  d  **  **
        1710: data = 8'b00111100; //  e   ****
        1711: data = 8'b00000000; //  f
          //    code x6b
        1712: data = 8'b00000000; //  0
        1713: data = 8'b00000000; //  1
        1714: data = 8'b11100000; //  2 ***
        1715: data = 8'b01100000; //  3  **
        1716: data = 8'b01100000; //  4  **
        1717: data = 8'b01100110; //  5  **  **
        1718: data = 8'b01101100; //  6  ** **
        1719: data = 8'b01111000; //  7  ****
        1720: data = 8'b01111000; //  8  ****
        1721: data = 8'b01101100; //  9  ** **
        1722: data = 8'b01100110; //  a  **  **
        1723: data = 8'b11100110; //  b ***  **
        1724: data = 8'b00000000; //  c
        1725: data = 8'b00000000; //  d
        1726: data = 8'b00000000; //  e
        1727: data = 8'b00000000; //  f
          //    code x6c
        1728: data = 8'b00000000; //  0
        1729: data = 8'b00000000; //  1
        1730: data = 8'b00111000; //  2   ***
        1731: data = 8'b00011000; //  3    **
        1732: data = 8'b00011000; //  4    **
        1733: data = 8'b00011000; //  5    **
        1734: data = 8'b00011000; //  6    **
        1735: data = 8'b00011000; //  7    **
        1736: data = 8'b00011000; //  8    **
        1737: data = 8'b00011000; //  9    **
        1738: data = 8'b00011000; //  a    **
        1739: data = 8'b00111100; //  b   ****
        1740: data = 8'b00000000; //  c
        1741: data = 8'b00000000; //  d
        1742: data = 8'b00000000; //  e
        1743: data = 8'b00000000; //  f
          //    code x6d
        1744: data = 8'b00000000; //  0
        1745: data = 8'b00000000; //  1
        1746: data = 8'b00000000; //  2
        1747: data = 8'b00000000; //  3
        1748: data = 8'b00000000; //  4
        1749: data = 8'b11100110; //  5 ***  **
        1750: data = 8'b11111111; //  6 ********
        1751: data = 8'b11011011; //  7 ** ** **
        1752: data = 8'b11011011; //  8 ** ** **
        1753: data = 8'b11011011; //  9 ** ** **
        1754: data = 8'b11011011; //  a ** ** **
        1755: data = 8'b11011011; //  b ** ** **
        1756: data = 8'b00000000; //  c
        1757: data = 8'b00000000; //  d
        1758: data = 8'b00000000; //  e
        1759: data = 8'b00000000; //  f
          //    code x6e
        1760: data = 8'b00000000; //  0
        1761: data = 8'b00000000; //  1
        1762: data = 8'b00000000; //  2
        1763: data = 8'b00000000; //  3
        1764: data = 8'b00000000; //  4
        1765: data = 8'b11011100; //  5 ** ***
        1766: data = 8'b01100110; //  6  **  **
        1767: data = 8'b01100110; //  7  **  **
        1768: data = 8'b01100110; //  8  **  **
        1769: data = 8'b01100110; //  9  **  **
        1770: data = 8'b01100110; //  a  **  **
        1771: data = 8'b01100110; //  b  **  **
        1772: data = 8'b00000000; //  c
        1773: data = 8'b00000000; //  d
        1774: data = 8'b00000000; //  e
        1775: data = 8'b00000000; //  f
          //    code x6f
        1776: data = 8'b00000000; //  0
        1777: data = 8'b00000000; //  1
        1778: data = 8'b00000000; //  2
        1779: data = 8'b00000000; //  3
        1780: data = 8'b00000000; //  4
        1781: data = 8'b01111100; //  5  *****
        1782: data = 8'b11000110; //  6 **   **
        1783: data = 8'b11000110; //  7 **   **
        1784: data = 8'b11000110; //  8 **   **
        1785: data = 8'b11000110; //  9 **   **
        1786: data = 8'b11000110; //  a **   **
        1787: data = 8'b01111100; //  b  *****
        1788: data = 8'b00000000; //  c
        1789: data = 8'b00000000; //  d
        1790: data = 8'b00000000; //  e
        1791: data = 8'b00000000; //  f
          //    code x70
        1792: data = 8'b00000000; //  0
        1793: data = 8'b00000000; //  1
        1794: data = 8'b00000000; //  2
        1795: data = 8'b00000000; //  3
        1796: data = 8'b00000000; //  4
        1797: data = 8'b11011100; //  5 ** ***
        1798: data = 8'b01100110; //  6  **  **
        1799: data = 8'b01100110; //  7  **  **
        1800: data = 8'b01100110; //  8  **  **
        1801: data = 8'b01100110; //  9  **  **
        1802: data = 8'b01100110; //  a  **  **
        1803: data = 8'b01111100; //  b  *****
        1804: data = 8'b01100000; //  c  **
        1805: data = 8'b01100000; //  d  **
        1806: data = 8'b11110000; //  e ****
        1807: data = 8'b00000000; //  f
          //    code x71
        1808: data = 8'b00000000; //  0
        1809: data = 8'b00000000; //  1
        1810: data = 8'b00000000; //  2
        1811: data = 8'b00000000; //  3
        1812: data = 8'b00000000; //  4
        1813: data = 8'b01110110; //  5  *** **
        1814: data = 8'b11001100; //  6 **  **
        1815: data = 8'b11001100; //  7 **  **
        1816: data = 8'b11001100; //  8 **  **
        1817: data = 8'b11001100; //  9 **  **
        1818: data = 8'b11001100; //  a **  **
        1819: data = 8'b01111100; //  b  *****
        1820: data = 8'b00001100; //  c     **
        1821: data = 8'b00001100; //  d     **
        1822: data = 8'b00011110; //  e    ****
        1823: data = 8'b00000000; //  f
          //    code x72
        1824: data = 8'b00000000; //  0
        1825: data = 8'b00000000; //  1
        1826: data = 8'b00000000; //  2
        1827: data = 8'b00000000; //  3
        1828: data = 8'b00000000; //  4
        1829: data = 8'b11011100; //  5 ** ***
        1830: data = 8'b01110110; //  6  *** **
        1831: data = 8'b01100110; //  7  **  **
        1832: data = 8'b01100000; //  8  **
        1833: data = 8'b01100000; //  9  **
        1834: data = 8'b01100000; //  a  **
        1835: data = 8'b11110000; //  b ****
        1836: data = 8'b00000000; //  c
        1837: data = 8'b00000000; //  d
        1838: data = 8'b00000000; //  e
        1839: data = 8'b00000000; //  f
          //    code x73
        1840: data = 8'b00000000; //  0
        1841: data = 8'b00000000; //  1
        1842: data = 8'b00000000; //  2
        1843: data = 8'b00000000; //  3
        1844: data = 8'b00000000; //  4
        1845: data = 8'b01111100; //  5  *****
        1846: data = 8'b11000110; //  6 **   **
        1847: data = 8'b01100000; //  7  **
        1848: data = 8'b00111000; //  8   ***
        1849: data = 8'b00001100; //  9     **
        1850: data = 8'b11000110; //  a **   **
        1851: data = 8'b01111100; //  b  *****
        1852: data = 8'b00000000; //  c
        1853: data = 8'b00000000; //  d
        1854: data = 8'b00000000; //  e
        1855: data = 8'b00000000; //  f
          //    code x74
        1856: data = 8'b00000000; //  0
        1857: data = 8'b00000000; //  1
        1858: data = 8'b00010000; //  2    *
        1859: data = 8'b00110000; //  3   **
        1860: data = 8'b00110000; //  4   **
        1861: data = 8'b11111100; //  5 ******
        1862: data = 8'b00110000; //  6   **
        1863: data = 8'b00110000; //  7   **
        1864: data = 8'b00110000; //  8   **
        1865: data = 8'b00110000; //  9   **
        1866: data = 8'b00110110; //  a   ** **
        1867: data = 8'b00011100; //  b    ***
        1868: data = 8'b00000000; //  c
        1869: data = 8'b00000000; //  d
        1870: data = 8'b00000000; //  e
        1871: data = 8'b00000000; //  f
          //    code x75
        1872: data = 8'b00000000; //  0
        1873: data = 8'b00000000; //  1
        1874: data = 8'b00000000; //  2
        1875: data = 8'b00000000; //  3
        1876: data = 8'b00000000; //  4
        1877: data = 8'b11001100; //  5 **  **
        1878: data = 8'b11001100; //  6 **  **
        1879: data = 8'b11001100; //  7 **  **
        1880: data = 8'b11001100; //  8 **  **
        1881: data = 8'b11001100; //  9 **  **
        1882: data = 8'b11001100; //  a **  **
        1883: data = 8'b01110110; //  b  *** **
        1884: data = 8'b00000000; //  c
        1885: data = 8'b00000000; //  d
        1886: data = 8'b00000000; //  e
        1887: data = 8'b00000000; //  f
          //    code x76
        1888: data = 8'b00000000; //  0
        1889: data = 8'b00000000; //  1
        1890: data = 8'b00000000; //  2
        1891: data = 8'b00000000; //  3
        1892: data = 8'b00000000; //  4
        1893: data = 8'b11000011; //  5 **    **
        1894: data = 8'b11000011; //  6 **    **
        1895: data = 8'b11000011; //  7 **    **
        1896: data = 8'b11000011; //  8 **    **
        1897: data = 8'b01100110; //  9  **  **
        1898: data = 8'b00111100; //  a   ****
        1899: data = 8'b00011000; //  b    **
        1900: data = 8'b00000000; //  c
        1901: data = 8'b00000000; //  d
        1902: data = 8'b00000000; //  e
        1903: data = 8'b00000000; //  f
          //    code x77
        1904: data = 8'b00000000; //  0
        1905: data = 8'b00000000; //  1
        1906: data = 8'b00000000; //  2
        1907: data = 8'b00000000; //  3
        1908: data = 8'b00000000; //  4
        1909: data = 8'b11000011; //  5 **    **
        1910: data = 8'b11000011; //  6 **    **
        1911: data = 8'b11000011; //  7 **    **
        1912: data = 8'b11011011; //  8 ** ** **
        1913: data = 8'b11011011; //  9 ** ** **
        1914: data = 8'b11111111; //  a ********
        1915: data = 8'b01100110; //  b  **  **
        1916: data = 8'b00000000; //  c
        1917: data = 8'b00000000; //  d
        1918: data = 8'b00000000; //  e
        1919: data = 8'b00000000; //  f
          //    code x78
        1920: data = 8'b00000000; //  0
        1921: data = 8'b00000000; //  1
        1922: data = 8'b00000000; //  2
        1923: data = 8'b00000000; //  3
        1924: data = 8'b00000000; //  4
        1925: data = 8'b11000011; //  5 **    **
        1926: data = 8'b01100110; //  6  **  **
        1927: data = 8'b00111100; //  7   ****
        1928: data = 8'b00011000; //  8    **
        1929: data = 8'b00111100; //  9   ****
        1930: data = 8'b01100110; //  a  **  **
        1931: data = 8'b11000011; //  b **    **
        1932: data = 8'b00000000; //  c
        1933: data = 8'b00000000; //  d
        1934: data = 8'b00000000; //  e
        1935: data = 8'b00000000; //  f
          //    code x79
        1936: data = 8'b00000000; //  0
        1937: data = 8'b00000000; //  1
        1938: data = 8'b00000000; //  2
        1939: data = 8'b00000000; //  3
        1940: data = 8'b00000000; //  4
        1941: data = 8'b11000110; //  5 **   **
        1942: data = 8'b11000110; //  6 **   **
        1943: data = 8'b11000110; //  7 **   **
        1944: data = 8'b11000110; //  8 **   **
        1945: data = 8'b11000110; //  9 **   **
        1946: data = 8'b11000110; //  a **   **
        1947: data = 8'b01111110; //  b  ******
        1948: data = 8'b00000110; //  c      **
        1949: data = 8'b00001100; //  d     **
        1950: data = 8'b11111000; //  e *****
        1951: data = 8'b00000000; //  f
          //    code x7a
        1952: data = 8'b00000000; //  0
        1953: data = 8'b00000000; //  1
        1954: data = 8'b00000000; //  2
        1955: data = 8'b00000000; //  3
        1956: data = 8'b00000000; //  4
        1957: data = 8'b11111110; //  5 *******
        1958: data = 8'b11001100; //  6 **  **
        1959: data = 8'b00011000; //  7    **
        1960: data = 8'b00110000; //  8   **
        1961: data = 8'b01100000; //  9  **
        1962: data = 8'b11000110; //  a **   **
        1963: data = 8'b11111110; //  b *******
        1964: data = 8'b00000000; //  c
        1965: data = 8'b00000000; //  d
        1966: data = 8'b00000000; //  e
        1967: data = 8'b00000000; //  f
          //    code x7b
        1968: data = 8'b00000000; //  0
        1969: data = 8'b00000000; //  1
        1970: data = 8'b00001110; //  2     ***
        1971: data = 8'b00011000; //  3    **
        1972: data = 8'b00011000; //  4    **
        1973: data = 8'b00011000; //  5    **
        1974: data = 8'b01110000; //  6  ***
        1975: data = 8'b00011000; //  7    **
        1976: data = 8'b00011000; //  8    **
        1977: data = 8'b00011000; //  9    **
        1978: data = 8'b00011000; //  a    **
        1979: data = 8'b00001110; //  b     ***
        1980: data = 8'b00000000; //  c
        1981: data = 8'b00000000; //  d
        1982: data = 8'b00000000; //  e
        1983: data = 8'b00000000; //  f
          //    code x7c
        1984: data = 8'b00000000; //  0
        1985: data = 8'b00000000; //  1
        1986: data = 8'b00011000; //  2    **
        1987: data = 8'b00011000; //  3    **
        1988: data = 8'b00011000; //  4    **
        1989: data = 8'b00011000; //  5    **
        1990: data = 8'b00000000; //  6
        1991: data = 8'b00011000; //  7    **
        1992: data = 8'b00011000; //  8    **
        1993: data = 8'b00011000; //  9    **
        1994: data = 8'b00011000; //  a    **
        1995: data = 8'b00011000; //  b    **
        1996: data = 8'b00000000; //  c
        1997: data = 8'b00000000; //  d
        1998: data = 8'b00000000; //  e
        1999: data = 8'b00000000; //  f
          //    code x7d
        2000: data = 8'b00000000; //  0
        2001: data = 8'b00000000; //  1
        2002: data = 8'b01110000; //  2  ***
        2003: data = 8'b00011000; //  3    **
        2004: data = 8'b00011000; //  4    **
        2005: data = 8'b00011000; //  5    **
        2006: data = 8'b00001110; //  6     ***
        2007: data = 8'b00011000; //  7    **
        2008: data = 8'b00011000; //  8    **
        2009: data = 8'b00011000; //  9    **
        2010: data = 8'b00011000; //  a    **
        2011: data = 8'b01110000; //  b  ***
        2012: data = 8'b00000000; //  c
        2013: data = 8'b00000000; //  d
        2014: data = 8'b00000000; //  e
        2015: data = 8'b00000000; //  f
          //    code x7e
        2016: data = 8'b00000000; //  0
        2017: data = 8'b00000000; //  1
        2018: data = 8'b01110110; //  2  *** **
        2019: data = 8'b11011100; //  3 ** ***
        2020: data = 8'b00000000; //  4
        2021: data = 8'b00000000; //  5
        2022: data = 8'b00000000; //  6
        2023: data = 8'b00000000; //  7
        2024: data = 8'b00000000; //  8
        2025: data = 8'b00000000; //  9
        2026: data = 8'b00000000; //  a
        2027: data = 8'b00000000; //  b
        2028: data = 8'b00000000; //  c
        2029: data = 8'b00000000; //  d
        2030: data = 8'b00000000; //  e
        2031: data = 8'b00000000; //  f
          //    code x7f
        2032: data = 8'b00000000; //  0
        2033: data = 8'b00000000; //  1
        2034: data = 8'b00000000; //  2
        2035: data = 8'b00000000; //  3
        2036: data = 8'b00010000; //  4    *
        2037: data = 8'b00111000; //  5   ***
        2038: data = 8'b01101100; //  6  ** **
        2039: data = 8'b11000110; //  7 **   **
        2040: data = 8'b11000110; //  8 **   **
        2041: data = 8'b11000110; //  9 **   **
        2042: data = 8'b11111110; //  a *******
        2043: data = 8'b00000000; //  b
        2044: data = 8'b00000000; //  c
        2045: data = 8'b00000000; //  d
        2046: data = 8'b00000000; //  e
        2047: data = 8'b00000000; //  f
    endcase
end
endmodule